# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2009, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *       NGLibraryCreator, v2009.07-HR28-2009-07-08 - build 0907160200        *
# *                                                                            *
# ******************************************************************************
# 
# 

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.0050 ;

LAYER metal1
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     0.3000     0.9000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.0650     0.0650     0.0650     0.0650     0.0650     0.0650     
      WIDTH 0.0900       0.0650     0.0900     0.0900     0.0900     0.0900     0.0900     
      WIDTH 0.2700       0.0650     0.0900     0.2700     0.2700     0.2700     0.2700     
      WIDTH 0.5000       0.0650     0.0900     0.2700     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.0650     0.0900     0.2700     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.0650     0.0900     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.07 ;
  PITCH 0.19 0.14 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.38 ;
  THICKNESS 0.13 ;
  HEIGHT 0.37 ;
  CAPACITANCE CPERSQDIST 7.71613e-05 ;
  EDGECAPACITANCE 3.86e-05 ;
END metal1

LAYER via1
  TYPE CUT ;
  SPACING 0.08 ;
  WIDTH 0.07 ;
  RESISTANCE 5 ;
END via1

LAYER metal2
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     0.3000     0.9000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.0700     0.0700     0.0700     0.0700     0.0700     0.0700     
      WIDTH 0.0900       0.0700     0.0900     0.0900     0.0900     0.0900     0.0900     
      WIDTH 0.2700       0.0700     0.0900     0.2700     0.2700     0.2700     0.2700     
      WIDTH 0.5000       0.0700     0.0900     0.2700     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.0700     0.0900     0.2700     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.0700     0.0900     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.07 ;
  PITCH 0.19 0.14 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.25 ;
  THICKNESS 0.14 ;
  HEIGHT 0.62 ;
  CAPACITANCE CPERSQDIST 4.08957e-05 ;
  EDGECAPACITANCE 2.04e-05 ;
END metal2

LAYER via2
  TYPE CUT ;
  SPACING 0.09 ;
  WIDTH 0.07 ;
  RESISTANCE 5 ;
END via2

LAYER metal3
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     0.3000     0.9000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.0700     0.0700     0.0700     0.0700     0.0700     0.0700     
      WIDTH 0.0900       0.0700     0.0900     0.0900     0.0900     0.0900     0.0900     
      WIDTH 0.2700       0.0700     0.0900     0.2700     0.2700     0.2700     0.2700     
      WIDTH 0.5000       0.0700     0.0900     0.2700     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.0700     0.0900     0.2700     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.0700     0.0900     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.07 ;
  PITCH 0.19 0.14 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.25 ;
  THICKNESS 0.14 ;
  HEIGHT 0.88 ;
  CAPACITANCE CPERSQDIST 2.7745e-05 ;
  EDGECAPACITANCE 1.39e-05 ;
END metal3

LAYER via3
  TYPE CUT ;
  SPACING 0.09 ;
  WIDTH 0.07 ;
  RESISTANCE 5 ;
END via3

LAYER metal4
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     0.9000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.1400     0.1400     0.1400     0.1400     0.1400     
      WIDTH 0.2700       0.1400     0.2700     0.2700     0.2700     0.2700     
      WIDTH 0.5000       0.1400     0.2700     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.1400     0.2700     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.1400     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.14 ;
  PITCH 0.28 0.28 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.21 ;
  THICKNESS 0.28 ;
  HEIGHT 1.14 ;
  CAPACITANCE CPERSQDIST 2.07429e-05 ;
  EDGECAPACITANCE 1.04e-05 ;
END metal4

LAYER via4
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
  RESISTANCE 3 ;
END via4

LAYER metal5
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     0.9000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.1400     0.1400     0.1400     0.1400     0.1400     
      WIDTH 0.2700       0.1400     0.2700     0.2700     0.2700     0.2700     
      WIDTH 0.5000       0.1400     0.2700     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.1400     0.2700     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.1400     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.14 ;
  PITCH 0.28 0.28 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.21 ;
  THICKNESS 0.28 ;
  HEIGHT 1.71 ;
  CAPACITANCE CPERSQDIST 1.3527e-05 ;
  EDGECAPACITANCE 6.76e-06 ;
END metal5

LAYER via5
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
  RESISTANCE 3 ;
END via5

LAYER metal6
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     0.9000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.1400     0.1400     0.1400     0.1400     0.1400     
      WIDTH 0.2700       0.1400     0.2700     0.2700     0.2700     0.2700     
      WIDTH 0.5000       0.1400     0.2700     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.1400     0.2700     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.1400     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.14 ;
  PITCH 0.28 0.28 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.21 ;
  THICKNESS 0.28 ;
  HEIGHT 2.28 ;
  CAPACITANCE CPERSQDIST 1.00359e-05 ;
  EDGECAPACITANCE 5.02e-06 ;
END metal6

LAYER via6
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
  RESISTANCE 3 ;
END via6

LAYER metal7
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.4000     0.4000     0.4000     0.4000     
      WIDTH 0.5000       0.4000     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.4000     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.4000     0.5000     0.9000     1.5000      ;
  WIDTH 0.4 ;
  PITCH 0.8 0.8 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.075 ;
  THICKNESS 0.8 ;
  HEIGHT 2.85 ;
  CAPACITANCE CPERSQDIST 7.97709e-06 ;
  EDGECAPACITANCE 3.99e-06 ;
END metal7

LAYER via7
  TYPE CUT ;
  SPACING 0.44 ;
  WIDTH 0.4 ;
  RESISTANCE 1 ;
END via7

LAYER metal8
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.4000     0.4000     0.4000     0.4000     
      WIDTH 0.5000       0.4000     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.4000     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.4000     0.5000     0.9000     1.5000      ;
  WIDTH 0.4 ;
  PITCH 0.8 0.8 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.075 ;
  THICKNESS 0.8 ;
  HEIGHT 4.47 ;
  CAPACITANCE CPERSQDIST 5.0391e-06 ;
  EDGECAPACITANCE 2.52e-06 ;
END metal8

LAYER via8
  TYPE CUT ;
  SPACING 0.44 ;
  WIDTH 0.4 ;
  RESISTANCE 1 ;
END via8

LAYER metal9
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     2.7000     4.0000     
      WIDTH 0.0000       0.8000     0.8000     0.8000     
      WIDTH 0.9000       0.8000     0.9000     0.9000     
      WIDTH 1.5000       0.8000     0.9000     1.5000      ;
  WIDTH 0.8 ;
  PITCH 1.6 1.6 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.03 ;
  THICKNESS 2 ;
  HEIGHT 6.09 ;
  CAPACITANCE CPERSQDIST 3.68273e-06 ;
  EDGECAPACITANCE 1.84e-06 ;
END metal9

LAYER via9
  TYPE CUT ;
  SPACING 0.88 ;
  WIDTH 0.8 ;
  RESISTANCE 0.5 ;
END via9

LAYER metal10
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     2.7000     4.0000     
      WIDTH 0.0000       0.8000     0.8000     0.8000     
      WIDTH 0.9000       0.8000     0.9000     0.9000     
      WIDTH 1.5000       0.8000     0.9000     1.5000      ;
  WIDTH 0.8 ;
  PITCH 1.6 1.6 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.03 ;
  THICKNESS 2 ;
  HEIGHT 10.09 ;
  CAPACITANCE CPERSQDIST 2.21236e-06 ;
  EDGECAPACITANCE 1.11e-06 ;
END metal10

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA via1_0 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via1_0

VIA via1_1 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via1_1

VIA via1_2 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via1_2

VIA via1_3 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal1 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER metal2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via1_3

VIA via1_4 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal1 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER metal2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via1_4

VIA via1_5 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal1 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER metal2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via1_5

VIA via1_6 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal1 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER metal2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via1_6

VIA via1_7 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal1 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER metal2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via1_7

VIA via1_8 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal1 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER metal2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via1_8

VIA via2_0 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via2_0

VIA via2_1 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via2_1

VIA via2_2 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via2_2

VIA via2_3 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER metal3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via2_3

VIA via2_4 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER metal3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via2_4

VIA via2_5 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via2_5

VIA via2_6 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER metal3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via2_6

VIA via2_7 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER metal3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via2_7

VIA via2_8 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via2_8

VIA via3_0 DEFAULT
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via3_0

VIA via3_1 DEFAULT
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via3_1

VIA via3_2 DEFAULT
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via3_2

VIA via4_0 DEFAULT
  LAYER via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via4_0

VIA via5_0 DEFAULT
  LAYER via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via5_0

VIA via6_0 DEFAULT
  LAYER via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END via6_0

VIA via7_0 DEFAULT
  LAYER via7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER metal7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER metal8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END via7_0

VIA via8_0 DEFAULT
  LAYER via8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER metal8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER metal9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
END via8_0

VIA via9_0 DEFAULT
  LAYER via9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER metal9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER metal10 ;
    RECT -0.4 -0.4 0.4 0.4 ;
END via9_0

VIARULE Via1Array-0 GENERATE
  LAYER metal1 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER metal2 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via1Array-0

VIARULE Via1Array-1 GENERATE
  LAYER metal1 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal2 ;
    ENCLOSURE 0 0.035 ;
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via1Array-1

VIARULE Via1Array-2 GENERATE
  LAYER metal1 ;
    ENCLOSURE 0.035 0 ;
  LAYER metal2 ;
    ENCLOSURE 0.035 0 ;
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via1Array-2

VIARULE Via1Array-3 GENERATE
  LAYER metal1 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal2 ;
    ENCLOSURE 0.035 0 ;
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via1Array-3

VIARULE Via1Array-4 GENERATE
  LAYER metal1 ;
    ENCLOSURE 0.035 0 ;
  LAYER metal2 ;
    ENCLOSURE 0 0.035 ;
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via1Array-4

VIARULE Via2Array-0 GENERATE
  LAYER metal2 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER metal3 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via2Array-0

VIARULE Via2Array-1 GENERATE
  LAYER metal2 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal3 ;
    ENCLOSURE 0 0.035 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via2Array-1

VIARULE Via2Array-2 GENERATE
  LAYER metal2 ;
    ENCLOSURE 0.035 0 ;
  LAYER metal3 ;
    ENCLOSURE 0.035 0 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via2Array-2

VIARULE Via2Array-3 GENERATE
  LAYER metal2 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal3 ;
    ENCLOSURE 0.035 0 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via2Array-3

VIARULE Via2Array-4 GENERATE
  LAYER metal2 ;
    ENCLOSURE 0.035 0 ;
  LAYER metal3 ;
    ENCLOSURE 0 0.035 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via2Array-4

VIARULE Via3Array-0 GENERATE
  LAYER metal3 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER metal4 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via3Array-0

VIARULE Via3Array-1 GENERATE
  LAYER metal3 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal4 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via3Array-1

VIARULE Via3Array-2 GENERATE
  LAYER metal3 ;
    ENCLOSURE 0.035 0 ;
  LAYER metal4 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via3Array-2

VIARULE Via4Array-0 GENERATE
  LAYER metal4 ;
    ENCLOSURE 0 0 ;
  LAYER metal5 ;
    ENCLOSURE 0 0 ;
  LAYER via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END Via4Array-0

VIARULE Via5Array-0 GENERATE
  LAYER metal5 ;
    ENCLOSURE 0 0 ;
  LAYER metal6 ;
    ENCLOSURE 0 0 ;
  LAYER via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END Via5Array-0

VIARULE Via6Array-0 GENERATE
  LAYER metal6 ;
    ENCLOSURE 0 0 ;
  LAYER metal7 ;
    ENCLOSURE 0.13 0.13 ;
  LAYER via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END Via6Array-0

VIARULE Via7Array-0 GENERATE
  LAYER metal7 ;
    ENCLOSURE 0 0 ;
  LAYER metal8 ;
    ENCLOSURE 0 0 ;
  LAYER via7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.84 BY 0.84 ;
END Via7Array-0

VIARULE Via8Array-0 GENERATE
  LAYER metal8 ;
    ENCLOSURE 0 0 ;
  LAYER metal9 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER via8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.84 BY 0.84 ;
END Via8Array-0

VIARULE Via9Array-0 GENERATE
  LAYER metal10 ;
    ENCLOSURE 0 0 ;
  LAYER metal9 ;
    ENCLOSURE 0 0 ;
  LAYER via9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
    SPACING 1.68 BY 1.68 ;
END Via9Array-0

SPACING
  SAMENET metal1 metal1 0.065 ;
  SAMENET metal2 metal2 0.07 ;
  SAMENET metal3 metal3 0.07 ;
  SAMENET metal4 metal4 0.14 ;
  SAMENET metal5 metal5 0.14 ;
  SAMENET metal6 metal6 0.14 ;
  SAMENET metal7 metal7 0.4 ;
  SAMENET metal8 metal8 0.4 ;
  SAMENET metal9 metal9 0.8 ;
  SAMENET metal10 metal10 0.8 ;
  SAMENET via1 via1 0.08 ;
  SAMENET via2 via2 0.09 ;
  SAMENET via3 via3 0.09 ;
  SAMENET via4 via4 0.16 ;
  SAMENET via5 via5 0.16 ;
  SAMENET via6 via6 0.16 ;
  SAMENET via7 via7 0.44 ;
  SAMENET via8 via8 0.44 ;
  SAMENET via9 via9 0.88 ;
  SAMENET via1 via2 0.0 STACK ;
  SAMENET via2 via3 0.0 STACK ;
  SAMENET via3 via4 0.0 STACK ;
  SAMENET via4 via5 0.0 STACK ;
  SAMENET via5 via6 0.0 STACK ;
  SAMENET via6 via7 0.0 STACK ;
  SAMENET via7 via8 0.0 STACK ;
  SAMENET via8 via9 0.0 STACK ;
END SPACING

SITE NCSU_FreePDK_45nm
  SYMMETRY y ;
  CLASS core ;
  SIZE 0.19 BY 1.4 ;
END NCSU_FreePDK_45nm

MACRO AND2_X1
  CLASS core ;
  FOREIGN AND2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.065 1.315 0.065 1.175 0.135 1.175 0.135 1.315 0.445 1.315 0.445 1.175 0.515 1.175 0.515 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.195 0.42 0.195 0.56 0.06 0.56  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.515 0.085 0.515 0.27 0.445 0.27 0.445 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.395 0.56 0.51 0.56 0.51 0.7 0.395 0.7  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.405 1.015 0.655 1.015 0.655 0.285 0.635 0.285 0.635 0.15 0.725 0.15 0.725 1.25 0.635 1.25 0.635 1.085 0.405 1.085  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.035 0.225 0.33 0.225 0.33 0.425 0.59 0.425 0.59 0.495 0.33 0.495 0.33 1.25 0.26 1.25 0.26 0.295 0.035 0.295  ;
  END
END AND2_X1

MACRO AND2_X2
  CLASS core ;
  FOREIGN AND2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.17 0.11 1.17 0.11 1.315 0.42 1.315 0.42 1.17 0.49 1.17 0.49 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.13 0.56 0.13 0.565 0.185 0.565 0.185 0.7 0.06 0.7  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.485 0.085 0.485 0.23 0.415 0.23 0.415 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.7 0.38 0.7 0.38 0.84 0.25 0.84  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.61 0.975 0.63 0.975 0.63 0.335 0.61 0.335 0.61 0.2 0.7 0.2 0.7 1.25 0.61 1.25  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.235 1.035 0.445 1.035 0.445 0.365 0.045 0.365 0.045 0.15 0.115 0.15 0.115 0.295 0.515 0.295 0.515 0.36 0.55 0.36 0.55 0.495 0.515 0.495 0.515 1.105 0.305 1.105 0.305 1.245 0.235 1.245  ;
  END
END AND2_X2

MACRO AND2_X4
  CLASS core ;
  FOREIGN AND2_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.065 1.315 0.065 1.175 0.135 1.175 0.135 1.315 0.44 1.315 0.44 1.175 0.51 1.175 0.51 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.13 0.56 0.13 0.705 0.185 0.705 0.185 0.84 0.06 0.84  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.51 0.085 0.51 0.195 0.44 0.195 0.44 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.7 0.43 0.7 0.43 0.84 0.25 0.84  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 0.205 0.7 0.205 0.7 0.985 0.63 0.985  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.26 1.04 0.495 1.04 0.495 0.33 0.035 0.33 0.035 0.15 0.17 0.15 0.17 0.26 0.565 0.26 0.565 1.11 0.33 1.11 0.33 1.25 0.26 1.25  ;
  END
END AND2_X4

MACRO AND3_X1
  CLASS core ;
  FOREIGN AND3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.225 1.315 0.225 1.175 0.295 1.175 0.295 1.315 0.605 1.315 0.605 1.175 0.675 1.175 0.675 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.7 0.595 0.7 0.595 0.84 0.44 0.84  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.495 0.215 0.495 0.215 0.63 0.13 0.63 0.13 0.7 0.06 0.7  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.675 0.085 0.675 0.27 0.605 0.27 0.605 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.7 0.28 0.7 0.28 0.51 0.405 0.51 0.405 0.645 0.35 0.645 0.35 0.84 0.25 0.84  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.8 1.115 0.82 1.115 0.82 0.285 0.8 0.285 0.8 0.15 0.89 0.15 0.89 1.25 0.8 1.25  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.045 1.04 0.66 1.04 0.66 0.41 0.045 0.41 0.045 0.22 0.11 0.22 0.11 0.34 0.755 0.34 0.755 0.475 0.73 0.475 0.73 1.11 0.485 1.11 0.485 1.25 0.415 1.25 0.415 1.11 0.115 1.11 0.115 1.25 0.045 1.25  ;
  END
END AND3_X1

MACRO AND3_X2
  CLASS core ;
  FOREIGN AND3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.225 1.315 0.225 1.17 0.295 1.17 0.295 1.315 0.605 1.315 0.605 1.17 0.675 1.17 0.675 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.405 0.67 0.595 0.67 0.595 0.805 0.405 0.805  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.185 0.42 0.185 0.56 0.06 0.56  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.675 0.085 0.675 0.195 0.605 0.195 0.605 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.42 0.38 0.42 0.38 0.56 0.25 0.56  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.8 0.975 0.82 0.975 0.82 0.3 0.8 0.3 0.8 0.165 0.89 0.165 0.89 1.25 0.8 1.25  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.045 1.035 0.66 1.035 0.66 0.355 0.045 0.355 0.045 0.155 0.115 0.155 0.115 0.285 0.73 0.285 0.73 0.565 0.74 0.565 0.74 0.7 0.73 0.7 0.73 1.105 0.49 1.105 0.49 1.245 0.42 1.245 0.42 1.105 0.115 1.105 0.115 1.245 0.045 1.245  ;
  END
END AND3_X2

MACRO AND3_X4
  CLASS core ;
  FOREIGN AND3_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.25 1.315 0.25 1.175 0.32 1.175 0.32 1.315 0.63 1.315 0.63 1.175 0.7 1.175 0.7 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.42 0.595 0.42 0.595 0.56 0.44 0.56  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.275 0.42 0.275 0.49 0.13 0.49 0.13 0.56 0.06 0.56  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.7 0.085 0.7 0.195 0.63 0.195 0.63 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.56 0.375 0.56 0.375 0.7 0.25 0.7  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.82 0.205 0.89 0.205 0.89 0.985 0.82 0.985  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.07 1 0.685 1 0.685 0.33 0.035 0.33 0.035 0.19 0.17 0.19 0.17 0.26 0.755 0.26 0.755 1.07 0.51 1.07 0.51 1.25 0.44 1.25 0.44 1.07 0.14 1.07 0.14 1.25 0.07 1.25  ;
  END
END AND3_X4

MACRO AND4_X1
  CLASS core ;
  FOREIGN AND4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.175 0.11 1.175 0.11 1.315 0.415 1.315 0.415 1.175 0.485 1.175 0.485 1.315 0.795 1.315 0.795 1.175 0.865 1.175 0.865 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.56 0.595 0.56 0.595 0.7 0.44 0.7  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.185 0.56 0.185 0.72 0.06 0.72  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.87 0.085 0.87 0.27 0.8 0.27 0.8 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.7 0.375 0.7 0.375 0.84 0.25 0.84  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.595 0.875 0.79 0.875 0.79 0.945 0.595 0.945  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.99 1.115 1.01 1.115 1.01 0.285 0.99 0.285 0.99 0.15 1.085 0.15 1.085 1.25 0.99 1.25  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.235 1.04 0.855 1.04 0.855 0.405 0.045 0.405 0.045 0.22 0.11 0.22 0.11 0.335 0.925 0.335 0.925 0.61 0.94 0.61 0.94 0.745 0.925 0.745 0.925 1.11 0.675 1.11 0.675 1.25 0.605 1.25 0.605 1.11 0.305 1.11 0.305 1.25 0.235 1.25  ;
  END
END AND4_X1

MACRO AND4_X2
  CLASS core ;
  FOREIGN AND4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.17 0.11 1.17 0.11 1.315 0.415 1.315 0.415 1.17 0.485 1.17 0.485 1.315 0.795 1.315 0.795 1.17 0.865 1.17 0.865 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.42 0.565 0.42 0.565 0.56 0.44 0.56  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.215 0.42 0.215 0.56 0.06 0.56  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.865 0.085 0.865 0.195 0.795 0.195 0.795 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.7 0.38 0.7 0.38 0.84 0.25 0.84  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 0.42 0.76 0.42 0.76 0.56 0.63 0.56  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.99 0.975 1.01 0.975 1.01 0.29 0.99 0.29 0.99 0.155 1.08 0.155 1.08 1.25 0.99 1.25  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.235 0.995 0.825 0.995 0.825 0.355 0.045 0.355 0.045 0.2 0.115 0.2 0.115 0.285 0.895 0.285 0.895 0.315 0.93 0.315 0.93 0.455 0.895 0.455 0.895 1.065 0.68 1.065 0.68 1.245 0.61 1.245 0.61 1.065 0.305 1.065 0.305 1.245 0.235 1.245  ;
  END
END AND4_X2

MACRO AND4_X4
  CLASS core ;
  FOREIGN AND4_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.175 0.11 1.175 0.11 1.315 0.415 1.315 0.415 1.175 0.485 1.175 0.485 1.315 0.795 1.315 0.795 1.175 0.865 1.175 0.865 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.42 0.565 0.42 0.565 0.56 0.44 0.56  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.13 0.42 0.13 0.585 0.19 0.585 0.19 0.72 0.06 0.72  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.865 0.085 0.865 0.195 0.795 0.195 0.795 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.42 0.325 0.42 0.325 0.585 0.38 0.585 0.38 0.72 0.255 0.72 0.255 0.56 0.25 0.56  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 0.42 0.7 0.42 0.7 0.555 0.755 0.555 0.755 0.69 0.63 0.69  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.99 0.71 1.01 0.71 1.01 0.45 0.99 0.45 0.99 0.175 1.08 0.175 1.08 0.985 0.99 0.985  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.235 1 0.825 1 0.825 0.355 0.045 0.355 0.045 0.2 0.115 0.2 0.115 0.285 0.895 0.285 0.895 0.475 0.93 0.475 0.93 0.61 0.895 0.61 0.895 1.07 0.675 1.07 0.675 1.25 0.605 1.25 0.605 1.07 0.305 1.07 0.305 1.25 0.235 1.25  ;
  END
END AND4_X4

MACRO ANTENNA_X1
  CLASS core ;
  FOREIGN ANTENNA_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.19 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.15 0.13 0.15 0.13 1.035 0.06 1.035  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.19 1.315 0.19 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.19 -0.085 0.19 0.085 0 0.085  ;
    END
  END VSS
END ANTENNA_X1

MACRO AOI211_X1
  CLASS core ;
  FOREIGN AOI211_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 0.84 0.845 0.84 0.845 0.98 0.63 0.98  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.82 1.315 0.82 1.165 0.89 1.165 0.89 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.705 0.085 0.705 0.27 0.635 0.27 0.635 0.085 0.135 0.085 0.135 0.23 0.065 0.23 0.065 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.555 0.56 0.7 0.56 0.7 0.7 0.555 0.7  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.22 0.625 0.42 0.625 0.42 0.15 0.51 0.15 0.51 0.35 0.82 0.35 0.82 0.15 0.89 0.15 0.89 0.42 0.49 0.42 0.49 0.695 0.29 0.695 0.29 1.015 0.355 1.015 0.355 1.085 0.22 1.085  ;
    END
  END ZN
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.24 0.42 0.24 0.56 0.06 0.56  ;
    END
  END C2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.365 0.795 0.545 0.795 0.545 0.945 0.365 0.945  ;
    END
  END C1
  OBS
      LAYER metal1 ;
        POLYGON 0.035 1.18 0.545 1.18 0.545 1.25 0.035 1.25  ;
  END
END AOI211_X1

MACRO AOI211_X2
  CLASS core ;
  FOREIGN AOI211_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.735 0.63 0.89 0.63 0.89 0.84 0.735 0.84  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.835 1.315 0.835 1.065 0.905 1.065 0.905 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.75 0.085 0.75 0.16 0.615 0.16 0.615 0.085 0.15 0.085 0.15 0.195 0.08 0.195 0.08 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.575 0.42 0.7 0.42 0.7 0.56 0.575 0.56  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.225 0.425 0.225 0.425 0.2 0.56 0.2 0.56 0.225 0.835 0.225 0.835 0.16 0.905 0.16 0.905 0.295 0.32 0.295 0.32 0.76 0.335 0.76 0.335 1.035 0.25 1.035  ;
    END
  END ZN
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.28 0.185 0.28 0.185 0.505 0.06 0.505  ;
    END
  END C2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.385 0.42 0.51 0.42 0.51 0.56 0.385 0.56  ;
    END
  END C1
  OBS
      LAYER metal1 ;
        POLYGON 0.085 0.945 0.155 0.945 0.155 1.15 0.46 1.15 0.46 0.945 0.53 0.945 0.53 1.22 0.085 1.22  ;
  END
END AOI211_X2

MACRO AOI211_X4
  CLASS core ;
  FOREIGN AOI211_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.71 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.065 0.42 1.27 0.42 1.27 0.575 1.065 0.575  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 1.145 1.315 1.145 1.24 1.28 1.24 1.28 1.315 1.71 1.315 1.71 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.71 -0.085 1.71 0.085 1.245 0.085 1.245 0.335 1.175 0.335 1.175 0.085 0.9 0.085 0.9 0.16 0.765 0.16 0.765 0.085 0.11 0.085 0.11 0.335 0.04 0.335 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.92 0.63 0.99 0.63 0.99 0.695 1.39 0.695 1.39 0.56 1.52 0.56 1.52 0.765 0.92 0.765  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2 0.905 0.785 0.905 0.785 0.35 0.39 0.35 0.39 0.28 1.09 0.28 1.09 0.35 0.89 0.35 0.89 0.42 0.855 0.42 0.855 0.975 0.2 0.975  ;
    END
  END ZN
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.15 0.63 0.22 0.63 0.22 0.77 0.63 0.77 0.63 0.63 0.72 0.63 0.72 0.84 0.15 0.84  ;
    END
  END C2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.315 0.56 0.51 0.56 0.51 0.7 0.315 0.7  ;
    END
  END C1
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.895 0.115 0.895 0.115 1.1 1.555 1.1 1.555 0.865 1.625 0.865 1.625 1.17 0.045 1.17  ;
  END
END AOI211_X4

MACRO AOI21_X1
  CLASS core ;
  FOREIGN AOI21_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.53 0.7 0.7 0.7 0.7 0.84 0.53 0.84  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.605 1.315 0.605 1.1 0.675 1.1 0.675 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.37 0.385 0.51 0.385 0.51 0.56 0.37 0.56  ;
    END
  END B1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.675 0.085 0.675 0.27 0.605 0.27 0.605 0.085 0.11 0.085 0.11 0.27 0.04 0.27 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.17 0.42 0.17 0.56 0.06 0.56  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.235 0.15 0.485 0.15 0.485 0.285 0.305 0.285 0.305 0.84 0.32 0.84 0.32 1.115 0.235 1.115  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.045 1.1 0.115 1.1 0.115 1.18 0.415 1.18 0.415 1.1 0.485 1.1 0.485 1.25 0.045 1.25  ;
  END
END AOI21_X1

MACRO AOI21_X2
  CLASS core ;
  FOREIGN AOI21_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.575 0.28 0.7 0.28 0.7 0.425 0.575 0.425  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.62 1.315 0.62 1.015 0.69 1.015 0.69 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.28 0.375 0.28 0.375 0.505 0.25 0.505  ;
    END
  END B1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.69 0.085 0.69 0.195 0.62 0.195 0.62 0.085 0.125 0.085 0.125 0.195 0.055 0.195 0.055 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.28 0.185 0.28 0.185 0.505 0.06 0.505  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.84 0.44 0.84 0.44 0.165 0.51 0.165 0.51 0.91 0.32 0.91 0.32 1.115 0.25 1.115  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.06 0.975 0.13 0.975 0.13 1.18 0.43 1.18 0.43 0.975 0.5 0.975 0.5 1.25 0.06 1.25  ;
  END
END AOI21_X2

MACRO AOI21_X4
  CLASS core ;
  FOREIGN AOI21_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.33 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.82 0.7 0.995 0.7 0.995 0.895 0.82 0.895  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.975 1.315 0.975 1.235 1.11 1.235 1.11 1.315 1.33 1.315 1.33 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.175 0.42 0.78 0.42 0.78 0.56 0.63 0.56 0.63 0.49 0.175 0.49  ;
    END
  END B1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.33 -0.085 1.33 0.085 1.075 0.085 1.075 0.335 1.005 0.335 1.005 0.085 0.54 0.085 0.54 0.16 0.405 0.16 0.405 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.56 0.51 0.56 0.51 0.7 0.44 0.7  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.04 0.245 0.92 0.245 0.92 0.315 0.11 0.315 0.11 0.84 0.13 0.84 0.13 0.915 0.73 0.915 0.73 0.985 0.04 0.985  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.065 1.08 1.195 1.08 1.195 0.92 1.265 0.92 1.265 1.15 0.135 1.15 0.135 1.22 0.065 1.22  ;
  END
END AOI21_X4

MACRO AOI221_X1
  CLASS core ;
  FOREIGN AOI221_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.405 0.595 0.565 0.595 0.565 0.73 0.495 0.73 0.495 0.665 0.405 0.665  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.23 1.315 0.23 1.16 0.3 1.16 0.3 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.42 0.325 0.42 0.325 0.73 0.405 0.73 0.405 0.865 0.255 0.865 0.255 0.56 0.25 0.56  ;
    END
  END B1
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.425 0.15 0.51 0.15 0.51 0.335 0.985 0.335 0.985 0.19 1.055 0.19 1.055 0.405 0.875 0.405 0.875 1.11 0.805 1.11 0.805 0.42 0.425 0.42  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.94 0.56 1.08 0.56 1.08 0.7 0.94 0.7  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.675 0.085 0.675 0.27 0.605 0.27 0.605 0.085 0.11 0.085 0.11 0.27 0.04 0.27 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.13 0.42 0.13 0.585 0.19 0.585 0.19 0.72 0.06 0.72  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 0.56 0.74 0.56 0.74 0.7 0.63 0.7  ;
    END
  END C2
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.975 0.485 0.975 0.485 1.25 0.415 1.25 0.415 1.045 0.115 1.045 0.115 1.25 0.045 1.25  ;
        POLYGON 0.615 0.975 0.685 0.975 0.685 1.18 0.985 1.18 0.985 0.975 1.055 0.975 1.055 1.25 0.615 1.25  ;
  END
END AOI221_X1

MACRO AOI221_X2
  CLASS core ;
  FOREIGN AOI221_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.56 0.595 0.56 0.595 0.7 0.44 0.7  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.225 1.315 0.225 1.205 0.295 1.205 0.295 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.63 0.375 0.63 0.375 0.84 0.25 0.84  ;
    END
  END B1
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.805 0.97 0.81 0.97 0.81 0.42 0.425 0.42 0.425 0.165 0.495 0.165 0.495 0.28 1.09 0.28 1.09 0.35 0.88 0.35 0.88 1.105 0.805 1.105  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.945 0.56 1.08 0.56 1.08 0.7 0.945 0.7  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.675 0.085 0.675 0.195 0.605 0.195 0.605 0.085 0.11 0.085 0.11 0.195 0.04 0.195 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.28 0.13 0.28 0.13 0.37 0.215 0.37 0.215 0.505 0.06 0.505  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.595 0.875 0.675 0.875 0.675 0.63 0.745 0.63 0.745 0.945 0.595 0.945  ;
    END
  END C2
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.77 0.115 0.77 0.115 1.045 0.52 1.045 0.52 1.115 0.045 1.115  ;
        POLYGON 0.58 1.17 1.09 1.17 1.09 1.24 0.58 1.24  ;
  END
END AOI221_X2

MACRO AOI221_X4
  CLASS core ;
  FOREIGN AOI221_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.09 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.96 0.63 1.03 0.63 1.03 0.705 1.905 0.705 1.905 0.56 2.03 0.56 2.03 0.775 0.96 0.775  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 1.225 1.315 1.225 1.205 1.665 1.205 1.665 1.315 2.09 1.315 2.09 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.54 0.28 1.65 0.28 1.65 0.42 1.61 0.42 1.61 0.505 1.54 0.505  ;
    END
  END B1
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.225 0.905 0.825 0.905 0.825 0.33 0.135 0.33 0.135 0.42 0.06 0.42 0.06 0.245 0.135 0.245 0.135 0.26 1.405 0.26 1.405 0.195 1.475 0.195 1.475 0.33 0.895 0.33 0.895 0.975 0.225 0.975  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.175 0.475 0.63 0.475 0.63 0.42 0.76 0.42 0.76 0.56 0.245 0.56 0.245 0.61 0.175 0.61  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.09 -0.085 2.09 0.085 1.855 0.085 1.855 0.195 1.785 0.195 1.785 0.085 1.1 0.085 1.1 0.195 1.03 0.195 1.03 0.085 0.51 0.085 0.51 0.195 0.44 0.195 0.44 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.105 0.57 1.71 0.57 1.71 0.505 1.765 0.505 1.765 0.42 1.84 0.42 1.84 0.64 1.105 0.64  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.545 0.63 0.7 0.63 0.7 0.84 0.545 0.84  ;
    END
  END C2
  OBS
      LAYER metal1 ;
        POLYGON 1 0.84 1.89 0.84 1.89 0.91 1 0.91  ;
        POLYGON 0.035 1.04 1.975 1.04 1.975 0.975 2.045 0.975 2.045 1.11 0.035 1.11  ;
  END
END AOI221_X4

MACRO AOI222_X1
  CLASS core ;
  FOREIGN AOI222_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.33 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.385 1.315 0.385 1.195 0.52 1.195 0.52 1.315 1.33 1.315 1.33 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 0.7 0.755 0.7 0.755 0.84 0.63 0.84  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.01 0.7 1.135 0.7 1.135 0.84 1.01 0.84  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.82 0.7 0.945 0.7 0.945 0.84 0.82 0.84  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.96 1.005 1.2 1.005 1.2 0.575 0.58 0.575 0.58 0.395 0.715 0.395 0.715 0.505 1.2 0.505 1.2 0.15 1.285 0.15 1.285 1.075 0.96 1.075  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.7 0.565 0.7 0.565 0.84 0.44 0.84  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.33 -0.085 1.33 0.085 0.93 0.085 0.93 0.195 0.795 0.195 0.795 0.085 0.335 0.085 0.335 0.405 0.2 0.405 0.2 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.7 0.185 0.7 0.185 0.84 0.06 0.84  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.7 0.375 0.7 0.375 0.84 0.25 0.84  ;
    END
  END C2
  OBS
      LAYER metal1 ;
        POLYGON 0.2 1.06 0.71 1.06 0.71 1.13 0.2 1.13  ;
        POLYGON 0.045 0.36 0.115 0.36 0.115 0.47 0.445 0.47 0.445 0.26 0.865 0.26 0.865 0.44 0.795 0.44 0.795 0.33 0.515 0.33 0.515 0.54 0.045 0.54  ;
        POLYGON 0.045 0.925 0.865 0.925 0.865 1.18 1.28 1.18 1.28 1.25 0.795 1.25 0.795 0.995 0.115 0.995 0.115 1.25 0.045 1.25  ;
  END
END AOI222_X1

MACRO AOI222_X2
  CLASS core ;
  FOREIGN AOI222_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.52 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.46 1.315 0.46 1.095 0.595 1.095 0.595 1.315 1.52 1.315 1.52 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.765 0.56 0.9 0.56 0.9 0.7 0.765 0.7  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.01 0.63 1.135 0.63 1.135 0.84 1.01 0.84  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.335 0.28 1.46 0.28 1.46 0.505 1.335 0.505  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.65 0.15 1.27 0.15 1.27 0.755 1.285 0.755 1.285 0.89 1.2 0.89 1.2 0.22 0.65 0.22  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6 0.42 0.7 0.42 0.7 0.56 0.6 0.56  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.52 -0.085 1.52 0.085 1.475 0.085 1.475 0.195 1.405 0.195 1.405 0.085 0.405 0.085 0.405 0.165 0.27 0.165 0.27 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.22 0.42 0.32 0.42 0.32 0.56 0.22 0.56  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.385 0.56 0.52 0.56 0.52 0.7 0.385 0.7  ;
    END
  END C2
  OBS
      LAYER metal1 ;
        POLYGON 0.27 0.785 0.78 0.785 0.78 0.855 0.27 0.855  ;
        POLYGON 0.08 0.285 0.97 0.285 0.97 0.355 0.08 0.355  ;
        POLYGON 0.115 0.755 0.185 0.755 0.185 0.96 1.405 0.96 1.405 0.755 1.475 0.755 1.475 1.03 1.05 1.03 1.05 1.245 0.915 1.245 0.915 1.03 0.115 1.03  ;
  END
END AOI222_X2

MACRO AOI222_X4
  CLASS core ;
  FOREIGN AOI222_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.66 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.22 1.315 0.22 1.1 0.355 1.1 0.355 1.315 0.605 1.315 0.605 1.1 0.74 1.1 0.74 1.315 2.66 1.315 2.66 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.2 0.56 1.27 0.56 1.27 0.7 1.2 0.7  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.88 0.525 1.95 0.525 1.95 0.625 2.34 0.625 2.34 0.56 2.52 0.56 2.52 0.7 1.88 0.7  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.085 0.42 2.22 0.42 2.22 0.56 2.085 0.56  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.805 0.79 2.625 0.79 2.625 0.86 1.72 0.86 1.72 0.35 0.415 0.35 0.415 0.28 2.625 0.28 2.625 0.35 1.84 0.35 1.84 0.42 1.805 0.42  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.405 0.455 0.545 0.455 0.545 0.525 0.405 0.525  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.66 -0.085 2.66 0.085 2.245 0.085 2.245 0.16 2.11 0.16 2.11 0.085 1.685 0.085 1.685 0.16 1.55 0.16 1.55 0.085 0.925 0.085 0.925 0.16 0.79 0.16 0.79 0.085 0.17 0.085 0.17 0.16 0.035 0.16 0.035 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.875 0.42 1.605 0.42 1.605 0.49 1.08 0.49 1.08 0.56 1.01 0.56 1.01 0.49 0.875 0.49  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.14 0.56 0.32 0.56 0.32 0.59 0.82 0.59 0.82 0.7 0.14 0.7  ;
    END
  END C2
  OBS
      LAYER metal1 ;
        POLYGON 0.07 0.77 0.14 0.77 0.14 0.85 1.65 0.85 1.65 1.015 1.58 1.015 1.58 0.92 0.07 0.92  ;
        POLYGON 0.985 1.08 2.435 1.08 2.435 1.15 0.985 1.15  ;
  END
END AOI222_X4

MACRO AOI22_X1
  CLASS core ;
  FOREIGN AOI22_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.24 1.315 0.24 1.1 0.31 1.1 0.31 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.28 0.375 0.28 0.375 0.725 0.305 0.725 0.305 0.42 0.25 0.42  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.575 0.28 0.7 0.28 0.7 0.42 0.575 0.42  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.88 0.085 0.88 0.23 0.81 0.23 0.81 0.085 0.125 0.085 0.125 0.23 0.055 0.23 0.055 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.13 0.42 0.13 0.485 0.23 0.485 0.23 0.62 0.06 0.62  ;
    END
  END B2
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.735 0.56 0.89 0.56 0.89 0.7 0.735 0.7  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.15 0.51 0.15 0.51 0.775 0.69 0.775 0.69 1.115 0.62 1.115 0.62 0.845 0.44 0.845  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.06 0.965 0.505 0.965 0.505 1.18 0.81 1.18 0.81 0.995 0.88 0.995 0.88 1.25 0.435 1.25 0.435 1.035 0.13 1.035 0.13 1.115 0.06 1.115  ;
  END
END AOI22_X1

MACRO AOI22_X2
  CLASS core ;
  FOREIGN AOI22_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.24 1.315 0.24 1.205 0.31 1.205 0.31 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.28 0.375 0.28 0.375 0.505 0.305 0.505 0.305 0.42 0.25 0.42  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.575 0.28 0.7 0.28 0.7 0.505 0.575 0.505  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.88 0.085 0.88 0.195 0.81 0.195 0.81 0.085 0.125 0.085 0.125 0.195 0.055 0.195 0.055 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.28 0.13 0.28 0.13 0.47 0.205 0.47 0.205 0.605 0.06 0.605  ;
    END
  END B2
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.765 0.28 0.89 0.28 0.89 0.505 0.765 0.505  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.245 0.51 0.245 0.51 0.92 0.725 0.92 0.725 0.99 0.44 0.99  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.06 1.055 0.88 1.055 0.88 1.19 0.81 1.19 0.81 1.125 0.13 1.125 0.13 1.19 0.06 1.19  ;
  END
END AOI22_X2

MACRO AOI22_X4
  CLASS core ;
  FOREIGN AOI22_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.71 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.195 1.315 0.195 1.24 0.33 1.24 0.33 1.315 0.575 1.315 0.575 1.24 0.71 1.24 0.71 1.315 1.71 1.315 1.71 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.215 0.595 0.44 0.595 0.44 0.665 0.215 0.665  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.2 0.56 1.43 0.56 1.43 0.63 1.27 0.63 1.27 0.7 1.2 0.7  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.71 -0.085 1.71 0.085 1.665 0.085 1.665 0.195 1.595 0.195 1.595 0.085 0.9 0.085 0.9 0.16 0.765 0.16 0.765 0.085 0.11 0.085 0.11 0.195 0.04 0.195 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.09 0.77 0.63 0.77 0.63 0.7 0.755 0.7 0.755 0.84 0.09 0.84  ;
    END
  END B2
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.955 0.765 1.39 0.765 1.39 0.7 1.62 0.7 1.62 0.84 0.955 0.84  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.89 0.92 1.51 0.92 1.51 0.99 0.82 0.99 0.82 0.35 0.39 0.35 0.39 0.28 1.32 0.28 1.32 0.35 0.89 0.35  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.045 1.005 0.115 1.005 0.115 1.07 1.595 1.07 1.595 1.005 1.665 1.005 1.665 1.14 0.045 1.14  ;
  END
END AOI22_X4

MACRO BUF_X1
  CLASS core ;
  FOREIGN BUF_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.42 0.15 0.51 0.15 0.51 1.25 0.42 1.25  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.22 0.56 0.22 0.7 0.06 0.7  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.195 1.315 0.195 1.21 0.33 1.21 0.33 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.33 0.085 0.33 0.235 0.195 0.235 0.195 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.045 1.075 0.285 1.075 0.285 0.37 0.045 0.37 0.045 0.15 0.115 0.15 0.115 0.3 0.355 0.3 0.355 1.145 0.115 1.145 0.115 1.25 0.045 1.25  ;
  END
END BUF_X1

MACRO BUF_X16
  CLASS core ;
  FOREIGN BUF_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.205 0.51 0.205 0.51 0.555 0.81 0.555 0.81 0.205 0.88 0.205 0.88 0.985 0.81 0.985 0.81 0.665 0.51 0.665 0.51 0.985 0.44 0.985  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.205 0.56 0.205 0.7 0.06 0.7  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.24 1.315 0.24 1.175 0.31 1.175 0.31 1.315 0.62 1.315 0.62 1.035 0.69 1.035 0.69 1.315 1 1.315 1 1.035 1.07 1.035 1.07 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 1.07 0.085 1.07 0.335 1 0.335 1 0.085 0.69 0.085 0.69 0.335 0.62 0.335 0.62 0.085 0.32 0.085 0.32 0.27 0.25 0.27 0.25 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.06 1.04 0.305 1.04 0.305 0.405 0.06 0.405 0.06 0.15 0.13 0.15 0.13 0.335 0.375 0.335 0.375 1.11 0.13 1.11 0.13 1.25 0.06 1.25  ;
  END
END BUF_X16

MACRO BUF_X2
  CLASS core ;
  FOREIGN BUF_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.42 0.975 0.44 0.975 0.44 0.3 0.42 0.3 0.42 0.165 0.51 0.165 0.51 1.25 0.42 1.25  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.215 0.56 0.215 0.7 0.06 0.7  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.225 1.315 0.225 1.17 0.295 1.17 0.295 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.3 0.085 0.3 0.285 0.23 0.285 0.23 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.045 1.035 0.28 1.035 0.28 0.495 0.045 0.495 0.045 0.165 0.115 0.165 0.115 0.425 0.375 0.425 0.375 0.56 0.35 0.56 0.35 1.105 0.115 1.105 0.115 1.245 0.045 1.245  ;
  END
END BUF_X2

MACRO BUF_X32
  CLASS core ;
  FOREIGN BUF_X32 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.71 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.425 0.255 0.495 0.255 0.495 0.57 0.8 0.57 0.8 0.255 0.87 0.255 0.87 0.57 1.175 0.57 1.175 0.255 1.245 0.255 1.245 0.57 1.555 0.57 1.555 0.255 1.625 0.255 1.625 0.94 1.555 0.94 1.555 0.685 1.245 0.685 1.245 0.94 1.175 0.94 1.175 0.685 0.87 0.685 0.87 0.94 0.8 0.94 0.8 0.685 0.495 0.685 0.495 0.94 0.425 0.94  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.19 0.56 0.19 0.7 0.06 0.7  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.225 1.315 0.225 1.175 0.295 1.175 0.295 1.315 0.605 1.315 0.605 1.065 0.675 1.065 0.675 1.315 0.995 1.315 0.995 1.065 1.065 1.065 1.065 1.315 1.365 1.315 1.365 1.065 1.435 1.065 1.435 1.315 1.71 1.315 1.71 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.71 -0.085 1.71 0.085 1.435 0.085 1.435 0.335 1.365 0.335 1.365 0.085 1.06 0.085 1.06 0.335 0.99 0.335 0.99 0.085 0.675 0.085 0.675 0.335 0.605 0.335 0.605 0.085 0.305 0.085 0.305 0.27 0.235 0.27 0.235 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.045 1.04 0.29 1.04 0.29 0.405 0.045 0.405 0.045 0.15 0.115 0.15 0.115 0.335 0.36 0.335 0.36 1.11 0.115 1.11 0.115 1.25 0.045 1.25  ;
  END
END BUF_X32

MACRO BUF_X4
  CLASS core ;
  FOREIGN BUF_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.435 0.74 0.44 0.74 0.44 0.555 0.435 0.555 0.435 0.28 0.51 0.28 0.51 1.015 0.435 1.015  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.205 0.56 0.205 0.7 0.06 0.7  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.24 1.315 0.24 1.175 0.31 1.175 0.31 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.31 0.085 0.31 0.27 0.24 0.27 0.24 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.06 1.04 0.27 1.04 0.27 0.405 0.06 0.405 0.06 0.15 0.13 0.15 0.13 0.335 0.34 0.335 0.34 0.58 0.375 0.58 0.375 0.715 0.34 0.715 0.34 1.11 0.13 1.11 0.13 1.25 0.06 1.25  ;
  END
END BUF_X4

MACRO BUF_X8
  CLASS core ;
  FOREIGN BUF_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.28 0.51 0.28 0.51 0.985 0.44 0.985  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.205 0.56 0.205 0.7 0.06 0.7  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.24 1.315 0.24 1.175 0.31 1.175 0.31 1.315 0.62 1.315 0.62 1.035 0.69 1.035 0.69 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.69 0.085 0.69 0.41 0.62 0.41 0.62 0.085 0.31 0.085 0.31 0.27 0.24 0.27 0.24 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.06 1.04 0.305 1.04 0.305 0.405 0.06 0.405 0.06 0.15 0.13 0.15 0.13 0.335 0.375 0.335 0.375 1.11 0.13 1.11 0.13 1.25 0.06 1.25  ;
  END
END BUF_X8

MACRO CLKBUF_X1
  CLASS core ;
  FOREIGN CLKBUF_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.15 0.52 0.15 0.52 1.25 0.44 1.25  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.24 0.56 0.24 0.7 0.06 0.7  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.235 1.315 0.235 1.21 0.37 1.21 0.37 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.37 0.085 0.37 0.235 0.235 0.235 0.235 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.035 1.075 0.305 1.075 0.305 0.37 0.035 0.37 0.035 0.185 0.17 0.185 0.17 0.3 0.375 0.3 0.375 1.145 0.17 1.145 0.17 1.215 0.035 1.215  ;
  END
END CLKBUF_X1

MACRO CLKBUF_X2
  CLASS core ;
  FOREIGN CLKBUF_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.42 0.975 0.44 0.975 0.44 0.3 0.42 0.3 0.42 0.165 0.51 0.165 0.51 1.25 0.42 1.25  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.19 0.56 0.19 0.7 0.06 0.7  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.23 1.315 0.23 1.17 0.3 1.17 0.3 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.3 0.085 0.3 0.285 0.23 0.285 0.23 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.045 1.035 0.255 1.035 0.255 0.495 0.045 0.495 0.045 0.165 0.115 0.165 0.115 0.425 0.375 0.425 0.375 0.59 0.325 0.59 0.325 1.105 0.115 1.105 0.115 1.245 0.045 1.245  ;
  END
END CLKBUF_X2

MACRO CLKBUF_X3
  CLASS core ;
  FOREIGN CLKBUF_X3 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.42 0.845 0.44 0.845 0.44 0.465 0.42 0.465 0.42 0.19 0.51 0.19 0.51 1.12 0.42 1.12  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.19 0.56 0.19 0.7 0.06 0.7  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.225 1.315 0.225 1.175 0.295 1.175 0.295 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.295 0.085 0.295 0.27 0.225 0.27 0.225 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.045 1.04 0.255 1.04 0.255 0.405 0.045 0.405 0.045 0.15 0.115 0.15 0.115 0.335 0.325 0.335 0.325 0.49 0.36 0.49 0.36 0.625 0.325 0.625 0.325 1.11 0.115 1.11 0.115 1.25 0.045 1.25  ;
  END
END CLKBUF_X3

MACRO CLKGATETST_X1
  CLASS core ;
  FOREIGN CLKGATETST_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.85 BY 1.4 ;
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.05 0.56 0.185 0.56 0.185 0.7 0.05 0.7  ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.385 1.315 0.385 1.21 0.52 1.21 0.52 1.315 1.145 1.315 1.145 1.21 1.28 1.21 1.28 1.315 1.7 1.315 1.7 1.115 1.835 1.115 1.835 1.315 2.045 1.315 2.045 1.115 2.18 1.115 2.18 1.315 2.425 1.315 2.425 1.115 2.56 1.115 2.56 1.315 2.85 1.315 2.85 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.85 -0.085 2.85 0.085 2.56 0.085 2.56 0.235 2.425 0.235 2.425 0.085 1.8 0.085 1.8 0.45 1.73 0.45 1.73 0.085 1.28 0.085 1.28 0.285 1.145 0.285 1.145 0.085 0.525 0.085 0.525 0.285 0.39 0.285 0.39 0.085 0.11 0.085 0.11 0.32 0.04 0.32 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN GCK
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.645 1.065 2.67 1.065 2.67 0.285 2.645 0.285 2.645 0.15 2.79 0.15 2.79 1.2 2.645 1.2  ;
    END
  END GCK
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.56 0.44 0.56 0.44 0.7 0.25 0.7  ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.15 0.56 2.225 0.56 2.225 0.7 2.15 0.7  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.8 0.505 0.8 0.505 0.42 0.2 0.42 0.2 0.325 0.335 0.325 0.335 0.35 0.575 0.35 0.575 0.87 0.115 0.87 0.115 1.075 0.045 1.075  ;
        POLYGON 0.74 1.18 1.01 1.18 1.01 1.075 1.47 1.075 1.47 1.145 1.08 1.145 1.08 1.25 0.67 1.25 0.67 0.155 1.01 0.155 1.01 0.35 1.365 0.35 1.365 0.285 1.435 0.285 1.435 0.42 1.01 0.42 1.01 0.55 0.94 0.55 0.94 0.225 0.74 0.225  ;
        POLYGON 0.805 0.29 0.875 0.29 0.875 0.755 1.485 0.755 1.485 0.89 0.875 0.89 0.875 1.115 0.805 1.115  ;
        POLYGON 1.065 0.615 1.55 0.615 1.55 0.42 1.62 0.42 1.62 1.02 1.55 1.02 1.55 0.685 1.065 0.685  ;
        POLYGON 1.875 0.15 2.01 0.15 2.01 0.22 1.99 0.22 1.99 1.02 1.92 1.02 1.92 0.22 1.875 0.22  ;
        POLYGON 2.27 0.885 2.29 0.885 2.29 0.375 2.08 0.375 2.08 0.24 2.36 0.24 2.36 0.725 2.605 0.725 2.605 0.86 2.36 0.86 2.36 1.02 2.27 1.02  ;
  END
END CLKGATETST_X1

MACRO CLKGATETST_X2
  CLASS core ;
  FOREIGN CLKGATETST_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.85 BY 1.4 ;
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.185 0.56 0.185 0.7 0.06 0.7  ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.385 1.315 0.385 1.07 0.52 1.07 0.52 1.315 1.145 1.315 1.145 1.21 1.28 1.21 1.28 1.315 1.7 1.315 1.7 1.035 1.835 1.035 1.835 1.315 2.045 1.315 2.045 0.975 2.18 0.975 2.18 1.315 2.425 1.315 2.425 1.115 2.56 1.115 2.56 1.315 2.85 1.315 2.85 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.85 -0.085 2.85 0.085 2.555 0.085 2.555 0.16 2.42 0.16 2.42 0.085 1.805 0.085 1.805 0.45 1.735 0.45 1.735 0.085 1.28 0.085 1.28 0.285 1.145 0.285 1.145 0.085 0.525 0.085 0.525 0.285 0.39 0.285 0.39 0.085 0.11 0.085 0.11 0.32 0.04 0.32 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN GCK
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.53 0.56 2.665 0.56 2.665 0.165 2.735 0.165 2.735 1.11 2.645 1.11 2.645 0.7 2.53 0.7  ;
    END
  END GCK
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.56 0.415 0.56 0.415 0.7 0.25 0.7  ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.15 0.56 2.225 0.56 2.225 0.7 2.15 0.7  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.8 0.5 0.8 0.5 0.42 0.2 0.42 0.2 0.325 0.335 0.325 0.335 0.35 0.57 0.35 0.57 0.87 0.115 0.87 0.115 1.075 0.045 1.075  ;
        POLYGON 0.73 1.18 1.01 1.18 1.01 1.075 1.47 1.075 1.47 1.145 1.08 1.145 1.08 1.25 0.66 1.25 0.66 0.155 1 0.155 1 0.35 1.365 0.35 1.365 0.285 1.435 0.285 1.435 0.42 1 0.42 1 0.55 0.93 0.55 0.93 0.225 0.73 0.225  ;
        POLYGON 0.795 0.29 0.865 0.29 0.865 0.68 1.48 0.68 1.48 0.815 0.865 0.815 0.865 1.115 0.795 1.115  ;
        POLYGON 1.065 0.545 1.545 0.545 1.545 0.42 1.615 0.42 1.615 1.08 1.545 1.08 1.545 0.615 1.065 0.615  ;
        POLYGON 1.87 0.15 2.005 0.15 2.005 0.22 1.99 0.22 1.99 0.94 1.92 0.94 1.92 0.22 1.87 0.22  ;
        POLYGON 2.27 0.885 2.29 0.885 2.29 0.39 2.08 0.39 2.08 0.165 2.15 0.165 2.15 0.32 2.6 0.32 2.6 0.39 2.36 0.39 2.36 1.02 2.27 1.02  ;
  END
END CLKGATETST_X2

MACRO CLKGATETST_X4
  CLASS core ;
  FOREIGN CLKGATETST_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.85 BY 1.4 ;
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.05 0.56 0.185 0.56 0.185 0.7 0.05 0.7  ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.385 1.315 0.385 0.93 0.52 0.93 0.52 1.315 1.145 1.315 1.145 1.07 1.28 1.07 1.28 1.315 1.695 1.315 1.695 1.085 1.83 1.085 1.83 1.315 2.075 1.315 2.075 0.94 2.145 0.94 2.145 1.315 2.415 1.315 2.415 0.975 2.55 0.975 2.55 1.315 2.85 1.315 2.85 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.85 -0.085 2.85 0.085 2.55 0.085 2.55 0.16 2.415 0.16 2.415 0.085 1.795 0.085 1.795 0.45 1.725 0.45 1.725 0.085 1.28 0.085 1.28 0.285 1.145 0.285 1.145 0.085 0.525 0.085 0.525 0.285 0.39 0.285 0.39 0.085 0.11 0.085 0.11 0.32 0.04 0.32 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN GCK
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.655 0.795 2.72 0.795 2.72 0.48 2.64 0.48 2.64 0.205 2.79 0.205 2.79 1.07 2.655 1.07  ;
    END
  END GCK
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.56 0.415 0.56 0.415 0.7 0.25 0.7  ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.15 0.42 2.22 0.42 2.22 0.68 2.15 0.68  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.765 0.5 0.765 0.5 0.425 0.2 0.425 0.2 0.325 0.335 0.325 0.335 0.355 0.57 0.355 0.57 0.835 0.115 0.835 0.115 1.04 0.045 1.04  ;
        POLYGON 0.74 1.18 1.01 1.18 1.01 0.935 1.47 0.935 1.47 1.005 1.08 1.005 1.08 1.25 0.67 1.25 0.67 0.155 1.01 0.155 1.01 0.35 1.335 0.35 1.335 0.325 1.47 0.325 1.47 0.42 1.01 0.42 1.01 0.55 0.94 0.55 0.94 0.225 0.74 0.225  ;
        POLYGON 0.805 0.29 0.875 0.29 0.875 0.71 1.48 0.71 1.48 0.845 0.875 0.845 0.875 1.115 0.805 1.115  ;
        POLYGON 1.1 0.485 1.545 0.485 1.545 0.42 1.615 0.42 1.615 1.14 1.545 1.14 1.545 0.62 1.1 0.62  ;
        POLYGON 1.875 0.15 2.01 0.15 2.01 0.22 1.99 0.22 1.99 0.99 1.92 0.99 1.92 0.22 1.875 0.22  ;
        POLYGON 2.265 0.795 2.285 0.795 2.285 0.355 2.075 0.355 2.075 0.22 2.355 0.22 2.355 0.53 2.595 0.53 2.595 0.6 2.355 0.6 2.355 0.93 2.265 0.93  ;
  END
END CLKGATETST_X4

MACRO CLKGATETST_X8
  CLASS core ;
  FOREIGN CLKGATETST_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 3.04 BY 1.4 ;
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.185 0.56 0.185 0.7 0.06 0.7  ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.385 1.315 0.385 1.205 0.52 1.205 0.52 1.315 1.145 1.315 1.145 1.065 1.28 1.065 1.28 1.315 1.675 1.315 1.675 1.005 1.81 1.005 1.81 1.315 2.02 1.315 2.02 0.975 2.155 0.975 2.155 1.315 2.395 1.315 2.395 0.84 2.53 0.84 2.53 1.315 2.805 1.315 2.805 0.945 2.875 0.945 2.875 1.315 3.04 1.315 3.04 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 3.04 -0.085 3.04 0.085 2.875 0.085 2.875 0.195 2.805 0.195 2.805 0.085 2.53 0.085 2.53 0.3 2.395 0.3 2.395 0.085 1.78 0.085 1.78 0.45 1.71 0.45 1.71 0.085 1.28 0.085 1.28 0.285 1.145 0.285 1.145 0.085 0.52 0.085 0.52 0.285 0.385 0.285 0.385 0.085 0.11 0.085 0.11 0.32 0.04 0.32 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN GCK
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.59 0.69 2.72 0.69 2.72 0.45 2.59 0.45 2.59 0.38 2.79 0.38 2.79 0.76 2.59 0.76  ;
    END
  END GCK
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.56 0.405 0.56 0.405 0.7 0.25 0.7  ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.77 0.545 1.85 0.545 1.85 0.7 1.77 0.7  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.765 0.5 0.765 0.5 0.485 0.235 0.485 0.235 0.29 0.305 0.29 0.305 0.415 0.57 0.415 0.57 0.835 0.115 0.835 0.115 1.04 0.045 1.04  ;
        POLYGON 0.73 1.175 1.01 1.175 1.01 0.93 1.435 0.93 1.435 1.25 1.365 1.25 1.365 1 1.08 1 1.08 1.245 0.66 1.245 0.66 0.155 1 0.155 1 0.35 1.365 0.35 1.365 0.285 1.435 0.285 1.435 0.42 1 0.42 1 0.55 0.93 0.55 0.93 0.225 0.73 0.225  ;
        POLYGON 0.795 0.29 0.865 0.29 0.865 0.62 1.485 0.62 1.485 0.755 0.87 0.755 0.87 1.11 0.795 1.11  ;
        POLYGON 1.525 0.81 1.55 0.81 1.55 0.555 1.065 0.555 1.065 0.485 1.525 0.485 1.525 0.42 1.62 0.42 1.62 0.945 1.525 0.945  ;
        POLYGON 1.9 0.775 1.915 0.775 1.915 0.45 1.9 0.45 1.9 0.22 1.85 0.22 1.85 0.15 1.985 0.15 1.985 0.91 1.9 0.91  ;
        POLYGON 2.055 0.15 2.235 0.15 2.235 0.555 2.615 0.555 2.615 0.625 2.34 0.625 2.34 0.76 2.165 0.76 2.165 0.285 2.055 0.285  ;
  END
END CLKGATETST_X8

MACRO CLKGATE_X1
  CLASS core ;
  FOREIGN CLKGATE_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.28 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.205 1.315 0.205 0.99 0.34 0.99 0.34 1.315 0.96 1.315 0.96 0.99 1.095 0.99 1.095 1.315 1.51 1.315 1.51 1.115 1.645 1.115 1.645 1.315 1.885 1.315 1.885 1.115 2.02 1.115 2.02 1.315 2.28 1.315 2.28 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.28 -0.085 2.28 0.085 2.04 0.085 2.04 0.2 1.905 0.2 1.905 0.085 1.645 0.085 1.645 0.41 1.51 0.41 1.51 0.085 1.095 0.085 1.095 0.285 0.96 0.285 0.96 0.085 0.335 0.085 0.335 0.285 0.2 0.285 0.2 0.085 0 0.085  ;
    END
  END VSS
  PIN GCK
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.09 1.095 2.15 1.095 2.15 0.22 2.105 0.22 2.105 0.15 2.24 0.15 2.24 1.165 2.09 1.165  ;
    END
  END GCK
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.82 0.42 0.955 0.42 0.955 0.56 0.82 0.56  ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.45 0.63 1.58 0.63 1.58 0.56 1.65 0.56 1.65 0.63 1.915 0.63 1.915 0.7 1.45 0.7  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.035 0.29 0.115 0.29 0.115 0.445 0.445 0.445 0.445 0.515 0.105 0.515 0.105 0.76 0.115 0.76 0.115 0.895 0.035 0.895  ;
        POLYGON 0.625 0.76 0.68 0.76 0.68 0.895 0.555 0.895 0.555 0.725 0.17 0.725 0.17 0.59 0.555 0.59 0.555 0.29 0.68 0.29 0.68 0.425 0.625 0.425  ;
        POLYGON 0.69 0.625 1.15 0.625 1.15 0.32 1.285 0.32 1.285 0.39 1.22 0.39 1.22 0.76 1.25 0.76 1.25 0.895 1.15 0.895 1.15 0.695 0.69 0.695  ;
        POLYGON 1.285 0.555 1.315 0.555 1.315 0.45 1.455 0.45 1.455 0.52 1.385 0.52 1.385 0.885 1.42 0.885 1.42 1.02 1.315 1.02 1.315 0.69 1.285 0.69  ;
        POLYGON 1.7 0.915 2.015 0.915 2.015 0.52 1.885 0.52 1.885 0.45 2.085 0.45 2.085 0.985 1.7 0.985  ;
  END
END CLKGATE_X1

MACRO CLKGATE_X2
  CLASS core ;
  FOREIGN CLKGATE_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.28 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.25 1.315 0.25 0.955 0.32 0.955 0.32 1.315 1 1.315 1 0.955 1.07 0.955 1.07 1.315 1.55 1.315 1.55 0.94 1.62 0.94 1.62 1.315 1.925 1.315 1.925 1.08 1.995 1.08 1.995 1.315 2.28 1.315 2.28 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.28 -0.085 2.28 0.085 2.015 0.085 2.015 0.365 1.945 0.365 1.945 0.085 1.605 0.085 1.605 0.195 1.535 0.195 1.535 0.085 1.07 0.085 1.07 0.32 1 0.32 1 0.085 0.31 0.085 0.31 0.32 0.24 0.32 0.24 0.085 0 0.085  ;
    END
  END VSS
  PIN GCK
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.135 0.975 2.14 0.975 2.14 0.525 1.925 0.525 1.925 0.455 2.135 0.455 2.135 0.335 2.21 0.335 2.21 1.11 2.135 1.11  ;
    END
  END GCK
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.82 0.28 0.89 0.28 0.89 0.375 0.965 0.375 0.965 0.55 0.82 0.55  ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.58 0.56 1.7 0.56 1.7 0.7 1.58 0.7  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.035 0.29 0.125 0.29 0.125 0.445 0.43 0.445 0.43 0.515 0.105 0.515 0.105 0.76 0.11 0.76 0.11 1.035 0.035 1.035  ;
        POLYGON 0.635 0.76 0.69 0.76 0.69 0.895 0.565 0.895 0.565 0.65 0.17 0.65 0.17 0.58 0.565 0.58 0.565 0.29 0.69 0.29 0.69 0.425 0.635 0.425  ;
        POLYGON 1.205 0.615 1.26 0.615 1.26 1.035 1.19 1.035 1.19 0.685 0.7 0.685 0.7 0.615 1.135 0.615 1.135 0.2 1.26 0.2 1.26 0.335 1.205 0.335  ;
        POLYGON 1.27 0.415 1.35 0.415 1.35 0.165 1.43 0.165 1.43 1.02 1.36 1.02 1.36 0.55 1.27 0.55  ;
        POLYGON 1.745 0.885 1.765 0.885 1.765 0.495 1.555 0.495 1.555 0.36 1.835 0.36 1.835 0.59 2.075 0.59 2.075 0.725 1.835 0.725 1.835 1.16 1.745 1.16  ;
  END
END CLKGATE_X2

MACRO CLKGATE_X4
  CLASS core ;
  FOREIGN CLKGATE_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.28 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.24 1.315 0.24 0.955 0.31 0.955 0.31 1.315 1 1.315 1 0.955 1.07 0.955 1.07 1.315 1.545 1.315 1.545 1.08 1.615 1.08 1.615 1.315 1.925 1.315 1.925 1.08 1.995 1.08 1.995 1.315 2.28 1.315 2.28 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.28 -0.085 2.28 0.085 1.995 0.085 1.995 0.455 1.925 0.455 1.925 0.085 1.6 0.085 1.6 0.195 1.53 0.195 1.53 0.085 1.07 0.085 1.07 0.32 1 0.32 1 0.085 0.31 0.085 0.31 0.32 0.24 0.32 0.24 0.085 0 0.085  ;
    END
  END VSS
  PIN GCK
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.925 0.875 2.12 0.875 2.12 0.205 2.19 0.205 2.19 1.07 2.12 1.07 2.12 0.945 1.925 0.945  ;
    END
  END GCK
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.82 0.28 0.89 0.28 0.89 0.375 0.965 0.375 0.965 0.55 0.895 0.55 0.895 0.505 0.82 0.505  ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.58 0.56 1.65 0.56 1.65 0.7 1.58 0.7  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.035 0.29 0.125 0.29 0.125 0.445 0.43 0.445 0.43 0.515 0.105 0.515 0.105 0.76 0.11 0.76 0.11 0.895 0.035 0.895  ;
        POLYGON 0.67 0.76 0.69 0.76 0.69 0.895 0.6 0.895 0.6 0.65 0.17 0.65 0.17 0.58 0.6 0.58 0.6 0.29 0.69 0.29 0.69 0.425 0.67 0.425  ;
        POLYGON 1.125 0.765 1.26 0.765 1.26 1.04 1.19 1.04 1.19 0.835 0.755 0.835 0.755 0.71 0.735 0.71 0.735 0.575 0.825 0.575 0.825 0.765 1.055 0.765 1.055 0.385 1.19 0.385 1.19 0.29 1.26 0.29 1.26 0.455 1.125 0.455  ;
        POLYGON 1.19 0.535 1.35 0.535 1.35 0.165 1.43 0.165 1.43 1.16 1.36 1.16 1.36 0.67 1.19 0.67  ;
        POLYGON 1.52 0.425 1.815 0.425 1.815 0.55 2.055 0.55 2.055 0.685 1.815 0.685 1.815 1.02 1.745 1.02 1.745 0.495 1.52 0.495  ;
  END
END CLKGATE_X4

MACRO CLKGATE_X8
  CLASS core ;
  FOREIGN CLKGATE_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.47 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.25 1.315 0.25 0.955 0.32 0.955 0.32 1.315 1.01 1.315 1.01 0.955 1.08 0.955 1.08 1.315 1.555 1.315 1.555 1.08 1.625 1.08 1.625 1.315 1.935 1.315 1.935 1.08 2.005 1.08 2.005 1.315 2.33 1.315 2.33 0.94 2.4 0.94 2.4 1.315 2.47 1.315 2.47 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.47 -0.085 2.47 0.085 2.4 0.085 2.4 0.335 2.33 0.335 2.33 0.085 2.025 0.085 2.025 0.46 1.955 0.46 1.955 0.085 1.61 0.085 1.61 0.195 1.54 0.195 1.54 0.085 1.08 0.085 1.08 0.32 1.01 0.32 1.01 0.085 0.32 0.085 0.32 0.32 0.25 0.32 0.25 0.085 0 0.085  ;
    END
  END VSS
  PIN GCK
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.15 0.205 2.22 0.205 2.22 1.07 2.15 1.07  ;
    END
  END GCK
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.82 0.42 0.975 0.42 0.975 0.56 0.82 0.56  ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.58 0.56 1.65 0.56 1.65 0.7 1.58 0.7  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.29 0.135 0.29 0.135 0.445 0.465 0.445 0.465 0.515 0.115 0.515 0.115 0.895 0.045 0.895  ;
        POLYGON 0.62 0.795 0.735 0.795 0.735 0.865 0.55 0.865 0.55 0.74 0.18 0.74 0.18 0.67 0.55 0.67 0.55 0.325 0.735 0.325 0.735 0.395 0.62 0.395  ;
        POLYGON 1.175 0.76 1.27 0.76 1.27 0.895 1.105 0.895 1.105 0.695 0.685 0.695 0.685 0.56 0.755 0.56 0.755 0.625 1.105 0.625 1.105 0.425 1.2 0.425 1.2 0.29 1.27 0.29 1.27 0.495 1.175 0.495  ;
        POLYGON 1.24 0.56 1.36 0.56 1.36 0.165 1.44 0.165 1.44 1.02 1.37 1.02 1.37 0.695 1.24 0.695  ;
        POLYGON 1.565 0.36 1.815 0.36 1.815 0.585 2.085 0.585 2.085 0.72 1.815 0.72 1.815 1.02 1.745 1.02 1.745 0.495 1.565 0.495  ;
  END
END CLKGATE_X8

MACRO DFFRS_X1
  CLASS core ;
  FOREIGN DFFRS_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 5.13 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.395 0.15 0.51 0.15 0.51 0.42 0.465 0.42 0.465 1.02 0.49 1.02 0.49 1.155 0.395 1.155  ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.71 0.635 0.78 0.635 0.78 0.7 1.48 0.7 1.48 0.84 1.39 0.84 1.39 0.77 0.71 0.77  ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.04 0.42 3.17 0.42 3.17 0.705 3.04 0.705  ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.235 1.315 0.235 1.08 0.305 1.08 0.305 1.315 0.575 1.315 0.575 1.08 0.645 1.08 0.645 1.315 0.95 1.315 0.95 1.08 1.02 1.08 1.02 1.315 1.3 1.315 1.3 1.155 1.37 1.155 1.37 1.315 1.835 1.315 1.835 0.95 1.905 0.95 1.905 1.315 2.61 1.315 2.61 1.08 2.68 1.08 2.68 1.315 3.15 1.315 3.15 1.08 3.22 1.08 3.22 1.315 3.84 1.315 3.84 1.06 3.975 1.06 3.975 1.315 4.63 1.315 4.63 1.025 4.7 1.025 4.7 1.315 5.01 1.315 5.01 1.205 5.08 1.205 5.08 1.315 5.13 1.315 5.13 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.05 0.15 0.13 0.15 0.13 1.155 0.05 1.155  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 5.13 -0.085 5.13 0.085 5.08 0.085 5.08 0.32 5.01 0.32 5.01 0.085 4.545 0.085 4.545 0.285 4.41 0.285 4.41 0.085 3.44 0.085 3.44 0.41 3.37 0.41 3.37 0.085 2.505 0.085 2.505 0.415 2.37 0.415 2.37 0.085 1.435 0.085 1.435 0.445 1.365 0.445 1.365 0.085 1.02 0.085 1.02 0.37 0.95 0.37 0.95 0.085 0.305 0.085 0.305 0.27 0.235 0.27 0.235 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 4.39 0.68 4.88 0.68 4.88 0.84 4.795 0.84 4.795 0.75 4.39 0.75  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.165 0.87 1.325 0.87 1.325 0.945 1.165 0.945  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.53 0.585 0.575 0.585 0.575 0.29 0.645 0.29 0.645 0.835 0.83 0.835 0.83 1.155 0.76 1.155 0.76 0.905 0.575 0.905 0.575 0.72 0.53 0.72  ;
        POLYGON 1.085 1.01 1.545 1.01 1.545 0.58 1.185 0.58 1.185 0.415 1.255 0.415 1.255 0.51 1.545 0.51 1.545 0.175 2.045 0.175 2.045 0.245 1.615 0.245 1.615 1.08 1.085 1.08  ;
        POLYGON 1.755 0.795 2.815 0.795 2.815 0.865 2.28 0.865 2.28 1.07 2.21 1.07 2.21 0.865 1.755 0.865 1.755 1.235 1.685 1.235 1.685 0.365 2.125 0.365 2.125 0.435 1.755 0.435  ;
        POLYGON 1.88 0.645 2.805 0.645 2.805 0.4 2.875 0.4 2.875 0.645 2.95 0.645 2.95 1.02 2.88 1.02 2.88 0.715 1.88 0.715  ;
        POLYGON 2.29 1.15 2.355 1.15 2.355 0.945 2.815 0.945 2.815 1.085 3.015 1.085 3.015 0.795 3.265 0.795 3.265 0.865 3.085 0.865 3.085 1.155 2.745 1.155 2.745 1.015 2.425 1.015 2.425 1.215 2.29 1.215  ;
        POLYGON 3.715 0.485 3.85 0.485 3.85 0.845 3.715 0.845  ;
        POLYGON 2.1 0.51 2.595 0.51 2.595 0.265 3.305 0.265 3.305 0.475 3.4 0.475 3.4 1.18 3.705 1.18 3.705 0.91 3.94 0.91 3.94 0.485 4.075 0.485 4.075 0.915 4.115 0.915 4.115 1.12 4.495 1.12 4.495 0.83 4.63 0.83 4.63 0.9 4.565 0.9 4.565 1.19 4.045 1.19 4.045 0.98 3.775 0.98 3.775 1.25 3.33 1.25 3.33 0.545 3.235 0.545 3.235 0.335 2.665 0.335 2.665 0.58 2.1 0.58  ;
        POLYGON 3.465 0.735 3.53 0.735 3.53 0.32 4.21 0.32 4.21 0.525 4.82 0.525 4.82 0.595 4.32 0.595 4.32 1.055 4.25 1.055 4.25 0.595 4.14 0.595 4.14 0.39 3.6 0.39 3.6 1.11 3.465 1.11  ;
        POLYGON 4.795 1.045 4.95 1.045 4.95 0.455 4.275 0.455 4.275 0.22 3.875 0.22 3.875 0.25 3.74 0.25 3.74 0.15 4.345 0.15 4.345 0.385 4.635 0.385 4.635 0.2 4.705 0.2 4.705 0.385 5.02 0.385 5.02 1.115 4.795 1.115  ;
  END
END DFFRS_X1

MACRO DFFRS_X2
  CLASS core ;
  FOREIGN DFFRS_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 5.13 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.035 0.21 0.13 0.21 0.13 0.45 0.11 0.45 0.11 0.945 0.035 0.945  ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.34 0.835 1.39 0.835 1.39 0.565 1.525 0.565 1.525 0.635 1.46 0.635 1.46 0.98 1.34 0.98  ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.04 0.585 3.205 0.585 3.205 0.69 3.04 0.69  ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.23 1.315 0.23 1.005 0.3 1.005 0.3 1.315 0.61 1.315 0.61 1.005 0.68 1.005 0.68 1.315 1.155 1.315 1.155 1.19 1.29 1.19 1.29 1.315 1.725 1.315 1.725 1.025 1.795 1.025 1.795 1.315 2.475 1.315 2.475 1.035 2.545 1.035 2.545 1.315 3.085 1.315 3.085 1.035 3.155 1.035 3.155 1.315 3.83 1.315 3.83 1.01 3.9 1.01 3.9 1.315 4.575 1.315 4.575 1.16 4.71 1.16 4.71 1.315 4.98 1.315 4.98 0.945 5.05 0.945 5.05 1.315 5.13 1.315 5.13 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.765 0.285 0.84 0.285 0.84 0.865 0.89 0.865 0.89 1.14 0.765 1.14  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 5.13 -0.085 5.13 0.085 4.595 0.085 4.595 0.285 4.46 0.285 4.46 0.085 3.405 0.085 3.405 0.36 3.055 0.36 3.055 0.085 2.395 0.085 2.395 0.41 2.26 0.41 2.26 0.085 1.395 0.085 1.395 0.365 1.26 0.365 1.26 0.085 1.015 0.085 1.015 0.32 0.945 0.32 0.945 0.085 0.295 0.085 0.295 0.395 0.225 0.395 0.225 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 4.24 0.645 4.375 0.645 4.375 0.87 4.24 0.87  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.135 0.835 1.19 0.835 1.19 0.565 1.325 0.565 1.325 0.635 1.27 0.635 1.27 0.98 1.135 0.98  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.175 0.65 0.605 0.65 0.605 0.315 0.675 0.315 0.675 0.72 0.485 0.72 0.485 1.08 0.415 1.08 0.415 0.785 0.175 0.785  ;
        POLYGON 1 0.43 1.1 0.43 1.1 0.365 1.17 0.365 1.17 0.43 1.475 0.43 1.475 0.175 1.88 0.175 1.88 0.245 1.545 0.245 1.545 0.5 1.07 0.5 1.07 1.095 1 1.095  ;
        POLYGON 1.68 0.885 2.135 0.885 2.135 0.75 2.75 0.75 2.75 0.82 2.205 0.82 2.205 1.11 2.07 1.11 2.07 0.955 1.635 0.955 1.635 1.095 1.565 1.095 1.565 0.885 1.61 0.885 1.61 0.36 1.98 0.36 1.98 0.43 1.68 0.43  ;
        POLYGON 1.765 0.615 2.63 0.615 2.63 0.42 2.7 0.42 2.7 0.615 2.885 0.615 2.885 0.975 2.815 0.975 2.815 0.685 1.9 0.685 1.9 0.78 1.765 0.78  ;
        POLYGON 2.15 1.18 2.34 1.18 2.34 0.9 2.68 0.9 2.68 1.04 2.95 1.04 2.95 0.765 3.205 0.765 3.205 0.835 3.02 0.835 3.02 1.11 2.61 1.11 2.61 0.97 2.41 0.97 2.41 1.25 2.15 1.25  ;
        POLYGON 3.675 0.44 3.81 0.44 3.81 0.81 3.675 0.81  ;
        POLYGON 2.025 0.48 2.475 0.48 2.475 0.285 2.835 0.285 2.835 0.44 3.34 0.44 3.34 1.18 3.665 1.18 3.665 0.875 3.965 0.875 3.965 0.51 3.875 0.51 3.875 0.44 4.035 0.44 4.035 1.165 4.44 1.165 4.44 0.715 4.565 0.715 4.565 0.85 4.51 0.85 4.51 1.235 3.965 1.235 3.965 0.945 3.735 0.945 3.735 1.25 3.27 1.25 3.27 0.51 2.765 0.51 2.765 0.355 2.545 0.355 2.545 0.55 2.025 0.55  ;
        POLYGON 3.425 1.025 3.49 1.025 3.49 0.3 4.17 0.3 4.17 0.49 4.945 0.49 4.945 0.655 4.875 0.655 4.875 0.56 4.17 0.56 4.17 0.94 4.32 0.94 4.32 1.005 4.1 1.005 4.1 0.37 3.56 0.37 3.56 1.095 3.425 1.095  ;
        POLYGON 4.8 0.72 5.01 0.72 5.01 0.42 4.325 0.42 4.325 0.235 3.71 0.235 3.71 0.165 4.395 0.165 4.395 0.35 4.985 0.35 4.985 0.2 5.08 0.2 5.08 0.79 4.87 0.79 4.87 1.065 4.8 1.065  ;
  END
END DFFRS_X2

MACRO DFFR_X1
  CLASS core ;
  FOREIGN DFFR_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 3.99 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.48 0.98 3.5 0.98 3.5 0.285 3.48 0.285 3.48 0.15 3.57 0.15 3.57 1.12 3.48 1.12  ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.99 0.49 3.1 0.49 3.1 0.42 3.17 0.42 3.17 0.56 2.99 0.56  ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.225 1.315 0.225 0.995 0.295 0.995 0.295 1.315 0.975 1.315 0.975 0.92 1.11 0.92 1.11 1.315 1.765 1.315 1.765 0.955 1.835 0.955 1.835 1.315 2.09 1.315 2.09 1.025 2.225 1.025 2.225 1.315 2.855 1.315 2.855 1.115 2.99 1.115 2.99 1.315 3.3 1.315 3.3 1.19 3.435 1.19 3.435 1.315 3.635 1.315 3.635 1.06 3.77 1.06 3.77 1.315 3.99 1.315 3.99 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.855 0.15 3.93 0.15 3.93 1.1 3.855 1.1  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 3.99 -0.085 3.99 0.085 3.77 0.085 3.77 0.235 3.635 0.235 3.635 0.085 3 0.085 3 0.36 2.865 0.36 2.865 0.085 2.225 0.085 2.225 0.355 2.09 0.355 2.09 0.085 1.87 0.085 1.87 0.325 1.735 0.325 1.735 0.085 0.925 0.085 0.925 0.375 0.79 0.375 0.79 0.085 0.33 0.085 0.33 0.16 0.195 0.16 0.195 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.69 0.58 1.875 0.58 1.875 0.665 1.69 0.665  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.175 0.56 0.32 0.56 0.32 0.7 0.175 0.7  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.04 0.165 0.11 0.165 0.11 0.345 0.59 0.345 0.59 0.48 0.11 0.48 0.11 0.935 0.04 0.935  ;
        POLYGON 0.435 0.63 0.655 0.63 0.655 0.27 0.4 0.27 0.4 0.2 0.725 0.2 0.725 0.63 1.22 0.63 1.22 0.7 0.505 0.7 0.505 1.115 0.435 1.115  ;
        POLYGON 1.375 0.755 2.3 0.755 2.3 0.825 1.49 0.825 1.49 0.97 1.355 0.97 1.355 0.85 0.685 0.85 0.685 1.25 0.36 1.25 0.36 1.18 0.615 1.18 0.615 0.78 1.3 0.78 1.3 0.325 1.49 0.325 1.49 0.395 1.375 0.395  ;
        POLYGON 1.9 0.89 2.365 0.89 2.365 0.525 1.955 0.525 1.955 0.465 1.625 0.465 1.625 0.64 1.44 0.64 1.44 0.57 1.555 0.57 1.555 0.395 2.025 0.395 2.025 0.455 2.435 0.455 2.435 0.89 2.655 0.89 2.655 1.05 2.585 1.05 2.585 0.96 2.035 0.96 2.035 0.985 1.9 0.985  ;
        POLYGON 2.475 1.115 2.72 1.115 2.72 0.355 2.47 0.355 2.47 0.285 2.79 0.285 2.79 0.64 3.265 0.64 3.265 0.775 2.79 0.775 2.79 1.185 2.475 1.185  ;
        POLYGON 2.855 0.915 2.925 0.915 2.925 0.98 3.335 0.98 3.335 0.415 3.24 0.415 3.24 0.21 3.405 0.21 3.405 0.64 3.435 0.64 3.435 0.775 3.405 0.775 3.405 1.05 3.23 1.05 3.23 1.2 3.095 1.2 3.095 1.05 2.855 1.05  ;
  END
END DFFR_X1

MACRO DFFR_X2
  CLASS core ;
  FOREIGN DFFR_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 3.99 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.45 1.04 3.725 1.04 3.725 0.42 3.67 0.42 3.67 0.32 3.45 0.32 3.45 0.2 3.585 0.2 3.585 0.25 3.795 0.25 3.795 1.11 3.45 1.11  ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.91 0.42 3.01 0.42 3.01 0.56 2.91 0.56  ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.175 1.315 0.175 1.03 0.33 1.03 0.33 1.315 0.915 1.315 0.915 0.99 1.05 0.99 1.05 1.315 1.72 1.315 1.72 0.955 1.79 0.955 1.79 1.315 2.03 1.315 2.03 1.065 2.165 1.065 2.165 1.315 2.85 1.315 2.85 1.065 2.985 1.065 2.985 1.315 3.25 1.315 3.25 1.01 3.385 1.01 3.385 1.315 3.635 1.315 3.635 1.24 3.77 1.24 3.77 1.315 3.99 1.315 3.99 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.86 0.165 3.93 0.165 3.93 1.145 3.86 1.145  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 3.99 -0.085 3.99 0.085 3.775 0.085 3.775 0.16 3.64 0.16 3.64 0.085 2.94 0.085 2.94 0.31 2.805 0.31 2.805 0.085 2.17 0.085 2.17 0.31 2.035 0.31 2.035 0.085 1.825 0.085 1.825 0.285 1.69 0.285 1.69 0.085 0.865 0.085 0.865 0.285 0.73 0.285 0.73 0.085 0.33 0.085 0.33 0.2 0.195 0.2 0.195 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.65 0.525 1.84 0.525 1.84 0.7 1.65 0.7  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.175 0.675 0.32 0.675 0.32 0.84 0.175 0.84  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.04 0.205 0.11 0.205 0.11 0.485 0.755 0.485 0.755 0.555 0.11 0.555 0.11 1.075 0.04 1.075  ;
        POLYGON 0.42 0.63 0.82 0.63 0.82 0.42 0.395 0.42 0.395 0.15 0.53 0.15 0.53 0.35 1.16 0.35 1.16 0.425 0.89 0.425 0.89 0.7 0.49 0.7 0.49 1.115 0.42 1.115  ;
        POLYGON 1.325 0.765 2.115 0.765 2.115 0.745 2.25 0.745 2.25 0.835 0.64 0.835 0.64 1.25 0.395 1.25 0.395 1.18 0.57 1.18 0.57 0.765 1.255 0.765 1.255 0.325 1.45 0.325 1.45 0.395 1.325 0.395  ;
        POLYGON 1.88 0.925 2.33 0.925 2.33 0.455 1.585 0.455 1.585 0.59 1.39 0.59 1.39 0.52 1.515 0.52 1.515 0.35 1.98 0.35 1.98 0.385 2.4 0.385 2.4 0.865 2.6 0.865 2.6 1 1.95 1 1.95 1.06 1.88 1.06  ;
        POLYGON 2.42 1.065 2.665 1.065 2.665 0.735 2.465 0.735 2.465 0.36 2.46 0.36 2.46 0.225 2.535 0.225 2.535 0.665 3.48 0.665 3.48 0.735 2.735 0.735 2.735 1.135 2.42 1.135  ;
        POLYGON 2.8 0.845 3.59 0.845 3.59 0.56 3.18 0.56 3.18 0.15 3.315 0.15 3.315 0.49 3.66 0.49 3.66 0.915 3.185 0.915 3.185 1.06 3.05 1.06 3.05 0.92 2.8 0.92  ;
  END
END DFFR_X2

MACRO DFFS_X1
  CLASS core ;
  FOREIGN DFFS_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 3.8 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.27 0.92 3.31 0.92 3.31 0.49 3.27 0.49 3.27 0.15 3.38 0.15 3.38 1.055 3.27 1.055  ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.72 0.84 2.9 0.84 2.9 0.98 2.72 0.98  ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.28 1.315 0.28 1.19 0.415 1.19 0.415 1.315 1.035 1.315 1.035 1.01 1.17 1.01 1.17 1.315 1.43 1.315 1.43 1.01 1.565 1.01 1.565 1.315 2.18 1.315 2.18 1.08 2.25 1.08 2.25 1.315 2.915 1.315 2.915 1.165 3.05 1.165 3.05 1.315 3.455 1.315 3.455 0.98 3.525 0.98 3.525 1.315 3.8 1.315 3.8 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.48 0.56 3.64 0.56 3.64 0.15 3.71 0.15 3.71 1.055 3.64 1.055 3.64 0.7 3.48 0.7  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 3.8 -0.085 3.8 0.085 3.53 0.085 3.53 0.27 3.46 0.27 3.46 0.085 2.98 0.085 2.98 0.41 2.845 0.41 2.845 0.085 2 0.085 2 0.41 1.865 0.41 1.865 0.085 1.145 0.085 1.145 0.405 1.075 0.405 1.075 0.085 0.35 0.085 0.35 0.28 0.215 0.28 0.215 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.41 0.4 0.41 0.4 0.835 0.46 0.835 0.46 0.97 0.33 0.97 0.33 0.56 0.25 0.56  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.58 0.42 1.65 0.42 1.65 0.675 1.58 0.675  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.065 0.285 0.135 0.285 0.135 1.035 0.525 1.035 0.525 0.87 0.67 0.87 0.67 0.435 0.74 0.435 0.74 0.94 0.595 0.94 0.595 1.105 0.065 1.105  ;
        POLYGON 0.66 1.005 0.805 1.005 0.805 0.37 0.6 0.37 0.6 0.3 0.875 0.3 0.875 0.665 1.31 0.665 1.31 0.6 1.38 0.6 1.38 0.735 0.875 0.735 0.875 1.075 0.66 1.075  ;
        POLYGON 0.965 0.81 1.445 0.81 1.445 0.285 1.515 0.285 1.515 0.945 0.965 0.945  ;
        POLYGON 1.62 0.81 1.715 0.81 1.715 0.22 1.285 0.22 1.285 0.54 0.94 0.54 0.94 0.235 0.535 0.235 0.535 0.74 0.465 0.74 0.465 0.165 1.01 0.165 1.01 0.47 1.215 0.47 1.215 0.15 1.785 0.15 1.785 0.795 2.065 0.795 2.065 0.22 2.495 0.22 2.495 0.29 2.135 0.29 2.135 0.88 1.62 0.88  ;
        POLYGON 1.775 0.945 2.2 0.945 2.2 0.48 2.275 0.48 2.275 0.36 2.41 0.36 2.41 0.48 3.07 0.48 3.07 0.615 3 0.615 3 0.55 2.27 0.55 2.27 0.945 2.63 0.945 2.63 1.2 2.56 1.2 2.56 1.015 1.775 1.015  ;
        POLYGON 2.335 0.685 3.135 0.685 3.135 0.415 3.045 0.415 3.045 0.345 3.205 0.345 3.205 0.65 3.245 0.65 3.245 0.79 3.205 0.79 3.205 1.25 3.135 1.25 3.135 0.755 2.405 0.755 2.405 0.88 2.335 0.88  ;
  END
END DFFS_X1

MACRO DFFS_X2
  CLASS core ;
  FOREIGN DFFS_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 3.8 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.285 0.965 3.43 0.965 3.43 0.56 3.285 0.56 3.285 0.165 3.36 0.165 3.36 0.49 3.505 0.49 3.505 1.03 3.355 1.03 3.355 1.25 3.285 1.25  ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.72 0.885 2.865 0.885 2.865 1.02 2.79 1.02 2.79 1.12 2.72 1.12  ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.225 1.315 0.225 1.155 0.295 1.155 0.295 1.315 1.015 1.315 1.015 1.115 1.15 1.115 1.15 1.315 1.395 1.315 1.395 0.935 1.53 0.935 1.53 1.315 2.145 1.315 2.145 1.06 2.28 1.06 2.28 1.315 2.94 1.315 2.94 1.025 3.01 1.025 3.01 1.315 3.47 1.315 3.47 1.17 3.54 1.17 3.54 1.315 3.8 1.315 3.8 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.66 0.975 3.67 0.975 3.67 0.3 3.66 0.3 3.66 0.165 3.74 0.165 3.74 1.25 3.66 1.25  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 3.8 -0.085 3.8 0.085 3.545 0.085 3.545 0.195 3.475 0.195 3.475 0.085 2.975 0.085 2.975 0.41 2.84 0.41 2.84 0.085 1.985 0.085 1.985 0.445 1.915 0.445 1.915 0.085 1.125 0.085 1.125 0.37 1.055 0.37 1.055 0.085 0.295 0.085 0.295 0.28 0.225 0.28 0.225 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.375 0.405 0.375 0.405 0.955 0.25 0.955  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.58 0.42 1.665 0.42 1.665 0.69 1.58 0.69  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.25 0.115 0.25 0.115 1.02 0.495 1.02 0.495 0.865 0.65 0.865 0.65 0.42 0.72 0.42 0.72 0.935 0.565 0.935 0.565 1.09 0.115 1.09 0.115 1.185 0.045 1.185  ;
        POLYGON 0.635 1 0.785 1 0.785 0.355 0.605 0.355 0.605 0.285 0.855 0.285 0.855 0.6 1.38 0.6 1.38 0.735 1.31 0.735 1.31 0.67 0.855 0.67 0.855 1.07 0.705 1.07 0.705 1.2 0.635 1.2  ;
        POLYGON 0.945 0.735 1.015 0.735 1.015 0.8 1.445 0.8 1.445 0.355 1.395 0.355 1.395 0.285 1.53 0.285 1.53 0.355 1.515 0.355 1.515 0.87 1.31 0.87 1.31 1.02 1.24 1.02 1.24 0.87 0.945 0.87  ;
        POLYGON 1.62 0.755 1.73 0.755 1.73 0.22 1.33 0.22 1.33 0.505 0.92 0.505 0.92 0.22 0.54 0.22 0.54 0.66 0.47 0.66 0.47 0.15 0.99 0.15 0.99 0.435 1.26 0.435 1.26 0.15 1.8 0.15 1.8 0.74 2.05 0.74 2.05 0.19 2.49 0.19 2.49 0.26 2.12 0.26 2.12 0.825 1.69 0.825 1.69 1.02 1.62 1.02  ;
        POLYGON 1.77 0.925 2.19 0.925 2.19 0.48 2.3 0.48 2.3 0.325 2.37 0.325 2.37 0.48 3.05 0.48 3.05 0.615 2.98 0.615 2.98 0.55 2.26 0.55 2.26 0.925 2.625 0.925 2.625 1.145 2.555 1.145 2.555 0.995 1.77 0.995  ;
        POLYGON 2.33 0.68 3.125 0.68 3.125 0.295 3.065 0.295 3.065 0.16 3.195 0.16 3.195 0.68 3.32 0.68 3.32 0.815 3.195 0.815 3.195 1.145 3.125 1.145 3.125 0.815 2.33 0.815  ;
  END
END DFFS_X2

MACRO DFF_X1
  CLASS core ;
  FOREIGN DFF_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 3.23 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.09 0.175 3.17 0.175 3.17 1.2 3.09 1.2  ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.2 1.315 0.2 1.1 0.335 1.1 0.335 1.315 0.955 1.315 0.955 1.115 1.09 1.115 1.09 1.315 1.55 1.315 1.55 1.115 1.685 1.115 1.685 1.315 2.31 1.315 2.31 1.115 2.445 1.115 2.445 1.315 2.86 1.315 2.86 1.115 2.995 1.115 2.995 1.315 3.23 1.315 3.23 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.71 0.175 2.795 0.175 2.795 1.155 2.71 1.155  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 3.23 -0.085 3.23 0.085 2.995 0.085 2.995 0.26 2.86 0.26 2.86 0.085 2.45 0.085 2.45 0.2 2.315 0.2 2.315 0.085 1.685 0.085 1.685 0.2 1.55 0.2 1.55 0.085 1.105 0.085 1.105 0.43 0.97 0.43 0.97 0.085 0.33 0.085 0.33 0.34 0.195 0.34 0.195 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.9 0.7 1.08 0.7 1.08 0.84 0.9 0.84  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.515 0.33 1.65 0.33 1.65 0.775 1.515 0.775  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.345 0.115 0.345 0.115 0.6 0.465 0.6 0.465 0.38 0.535 0.38 0.535 0.83 0.465 0.83 0.465 0.69 0.115 0.69 0.115 1.185 0.045 1.185  ;
        POLYGON 0.615 1.05 0.63 1.05 0.63 0.255 0.7 0.255 0.7 0.905 1.18 0.905 1.18 0.975 0.7 0.975 0.7 1.185 0.615 1.185  ;
        POLYGON 0.765 0.545 1.195 0.545 1.195 0.345 1.315 0.345 1.315 1.2 1.245 1.2 1.245 0.615 0.835 0.615 0.835 0.68 0.765 0.68  ;
        POLYGON 1.45 0.84 1.81 0.84 1.81 0.29 2.105 0.29 2.105 0.425 1.925 0.425 1.925 0.91 1.465 0.91 1.465 1.02 1.38 1.02 1.38 0.22 1.195 0.22 1.195 0.15 1.46 0.15 1.46 0.285 1.45 0.285  ;
        POLYGON 1.935 1.115 2.17 1.115 2.17 0.22 1.93 0.22 1.93 0.15 2.24 0.15 2.24 0.69 2.47 0.69 2.47 0.825 2.24 0.825 2.24 1.185 1.935 1.185  ;
        POLYGON 2.305 0.42 2.535 0.42 2.535 0.15 2.605 0.15 2.605 0.42 2.645 0.42 2.645 0.555 2.605 0.555 2.605 1.2 2.535 1.2 2.535 0.555 2.305 0.555  ;
  END
END DFF_X1

MACRO DFF_X2
  CLASS core ;
  FOREIGN DFF_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 3.23 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.91 0.42 3.07 0.42 3.07 0.165 3.14 0.165 3.14 1.16 3.07 1.16 3.07 0.56 2.91 0.56  ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.215 1.315 0.215 1.04 0.35 1.04 0.35 1.315 0.98 1.315 0.98 1.115 1.115 1.115 1.115 1.315 1.535 1.315 1.535 1.115 1.67 1.115 1.67 1.315 2.305 1.315 2.305 0.935 2.44 0.935 2.44 1.315 2.855 1.315 2.855 0.975 2.99 0.975 2.99 1.315 3.23 1.315 3.23 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.7 0.165 2.79 0.165 2.79 1.16 2.7 1.16  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 3.23 -0.085 3.23 0.085 2.99 0.085 2.99 0.16 2.855 0.16 2.855 0.085 2.44 0.085 2.44 0.2 2.305 0.2 2.305 0.085 1.675 0.085 1.675 0.2 1.54 0.2 1.54 0.085 1.11 0.085 1.11 0.375 0.975 0.375 0.975 0.085 0.35 0.085 0.35 0.365 0.215 0.365 0.215 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.87 0.705 1.115 0.705 1.115 0.805 0.87 0.805  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.515 0.33 1.65 0.33 1.65 0.895 1.515 0.895  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.065 0.295 0.135 0.295 0.135 0.585 0.615 0.585 0.615 0.72 0.135 0.72 0.135 1.035 0.065 1.035  ;
        POLYGON 0.6 1.02 0.695 1.02 0.695 0.385 0.6 0.385 0.6 0.315 0.765 0.315 0.765 0.5 1.18 0.5 1.18 0.635 0.765 0.635 0.765 1.09 0.6 1.09  ;
        POLYGON 0.325 0.825 0.485 0.825 0.485 1.175 0.84 1.175 0.84 0.96 1.245 0.96 1.245 0.425 1.2 0.425 1.2 0.29 1.315 0.29 1.315 1.2 1.2 1.2 1.2 1.03 0.91 1.03 0.91 1.245 0.415 1.245 0.415 0.895 0.325 0.895  ;
        POLYGON 1.21 0.15 1.45 0.15 1.45 0.96 1.82 0.96 1.82 0.29 2.095 0.29 2.095 0.36 1.89 0.36 1.89 1.03 1.38 1.03 1.38 0.22 1.21 0.22  ;
        POLYGON 1.955 0.685 2.16 0.685 2.16 0.22 1.92 0.22 1.92 0.15 2.23 0.15 2.23 0.64 2.485 0.64 2.485 0.78 2.025 0.78 2.025 1.02 1.955 1.02  ;
        POLYGON 2.525 0.885 2.55 0.885 2.55 0.555 2.295 0.555 2.295 0.42 2.52 0.42 2.52 0.29 2.635 0.29 2.635 1.02 2.525 1.02  ;
  END
END DFF_X2

MACRO DLH_X1
  CLASS core ;
  FOREIGN DLH_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.09 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.22 1.315 0.22 1.1 0.355 1.1 0.355 1.315 0.57 1.315 0.57 1.1 0.705 1.1 0.705 1.315 1.325 1.315 1.325 1.1 1.46 1.1 1.46 1.315 1.7 1.315 1.7 1.21 1.835 1.21 1.835 1.315 2.09 1.315 2.09 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.77 0.56 1.915 0.56 1.915 0.15 1.985 0.15 1.985 1.25 1.915 1.25 1.915 0.7 1.77 0.7  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.09 -0.085 2.09 0.085 1.835 0.085 1.835 0.235 1.7 0.235 1.7 0.085 1.46 0.085 1.46 0.16 1.325 0.16 1.325 0.085 0.705 0.085 0.705 0.16 0.57 0.16 0.57 0.085 0.36 0.085 0.36 0.185 0.225 0.185 0.225 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.685 0.28 0.89 0.28 0.89 0.42 0.755 0.42 0.755 0.9 0.685 0.9  ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.215 0.42 0.215 0.56 0.06 0.56  ;
    END
  END G
  OBS
      LAYER metal1 ;
        POLYGON 0.07 0.65 0.28 0.65 0.28 0.32 0.035 0.32 0.035 0.225 0.17 0.225 0.17 0.25 0.35 0.25 0.35 0.65 0.465 0.65 0.465 0.72 0.14 0.72 0.14 1.195 0.07 1.195  ;
        POLYGON 0.41 0.955 0.545 0.955 0.545 0.295 0.415 0.295 0.415 0.225 0.615 0.225 0.615 0.965 0.85 0.965 0.85 0.825 1.165 0.825 1.165 0.895 0.92 0.895 0.92 1.035 0.41 1.035  ;
        POLYGON 0.985 0.96 1.23 0.96 1.23 0.525 0.985 0.525 0.985 0.165 1.055 0.165 1.055 0.455 1.48 0.455 1.48 0.59 1.3 0.59 1.3 1.03 1.055 1.03 1.055 1.235 0.985 1.235  ;
        POLYGON 1.22 0.275 1.615 0.275 1.615 1.165 1.545 1.165 1.545 0.39 1.22 0.39  ;
  END
END DLH_X1

MACRO DLH_X2
  CLASS core ;
  FOREIGN DLH_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.09 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.245 1.315 0.245 1.24 0.38 1.24 0.38 1.315 0.585 1.315 0.585 1.24 0.72 1.24 0.72 1.315 1.34 1.315 1.34 1.1 1.475 1.1 1.475 1.315 1.74 1.315 1.74 1.15 1.875 1.15 1.875 1.315 2.09 1.315 2.09 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.96 0.215 2.03 0.215 2.03 1.195 1.96 1.195  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.09 -0.085 2.09 0.085 1.875 0.085 1.875 0.21 1.74 0.21 1.74 0.085 1.475 0.085 1.475 0.16 1.34 0.16 1.34 0.085 0.685 0.085 0.685 0.195 0.615 0.195 0.615 0.085 0.38 0.085 0.38 0.16 0.245 0.16 0.245 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 0.7 0.695 0.7 0.695 0.29 0.765 0.29 0.765 0.895 0.63 0.895  ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.24 0.56 0.24 0.7 0.06 0.7  ;
    END
  END G
  OBS
      LAYER metal1 ;
        POLYGON 0.055 0.95 0.33 0.95 0.33 0.385 0.055 0.385 0.055 0.2 0.19 0.2 0.19 0.315 0.4 0.315 0.4 1.02 0.19 1.02 0.19 1.16 0.055 1.16  ;
        POLYGON 0.535 1.015 0.83 1.015 0.83 0.83 1.18 0.83 1.18 0.9 0.9 0.9 0.9 1.085 0.535 1.085 0.535 1.195 0.465 1.195 0.465 0.165 0.535 0.165 0.535 0.44 0.595 0.44 0.595 0.575 0.535 0.575  ;
        POLYGON 1 0.965 1.245 0.965 1.245 0.525 1 0.525 1 0.165 1.07 0.165 1.07 0.455 1.52 0.455 1.52 0.59 1.315 0.59 1.315 1.035 1.07 1.035 1.07 1.24 1 1.24  ;
        POLYGON 1.235 0.25 1.685 0.25 1.685 0.32 1.655 0.32 1.655 1.195 1.585 1.195 1.585 0.39 1.235 0.39  ;
  END
END DLH_X2

MACRO DLL_X1
  CLASS core ;
  FOREIGN DLL_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.9 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.195 1.315 0.195 1.065 0.33 1.065 0.33 1.315 0.54 1.315 0.54 1.115 0.675 1.115 0.675 1.315 1.295 1.315 1.295 1.115 1.43 1.115 1.43 1.315 1.55 1.315 1.55 0.945 1.685 0.945 1.685 1.315 1.9 1.315 1.9 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.765 0.37 1.84 0.37 1.84 1.03 1.765 1.03  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.9 -0.085 1.9 0.085 1.69 0.085 1.69 0.46 1.555 0.46 1.555 0.085 1.445 0.085 1.445 0.285 1.31 0.285 1.31 0.085 0.64 0.085 0.64 0.32 0.57 0.32 0.57 0.085 0.33 0.085 0.33 0.21 0.195 0.21 0.195 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 0.7 0.78 0.7 0.78 0.84 0.63 0.84  ;
    END
  END D
  PIN GN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.22 0.56 0.22 0.7 0.06 0.7  ;
    END
  END GN
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.825 0.285 0.825 0.285 0.35 0.045 0.35 0.045 0.215 0.115 0.215 0.115 0.28 0.355 0.28 0.355 0.895 0.115 0.895 0.115 1.11 0.045 1.11  ;
        POLYGON 0.385 0.955 0.42 0.955 0.42 0.215 0.49 0.215 0.49 0.955 0.845 0.955 0.845 0.61 0.915 0.61 0.915 1.025 0.385 1.025  ;
        POLYGON 0.955 1.08 0.98 1.08 0.98 0.425 0.95 0.425 0.95 0.29 1.05 0.29 1.05 0.61 1.335 0.61 1.335 0.745 1.05 0.745 1.05 1.215 0.955 1.215  ;
        POLYGON 1.19 0.97 1.4 0.97 1.4 0.455 1.205 0.455 1.205 0.36 1.48 0.36 1.48 1.04 1.19 1.04  ;
  END
END DLL_X1

MACRO DLL_X2
  CLASS core ;
  FOREIGN DLL_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.9 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.195 1.315 0.195 1.02 0.33 1.02 0.33 1.315 0.575 1.315 0.575 1.08 0.645 1.08 0.645 1.315 1.3 1.315 1.3 1.115 1.435 1.115 1.435 1.315 1.6 1.315 1.6 0.91 1.67 0.91 1.67 1.315 1.9 1.315 1.9 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.77 0.28 1.85 0.28 1.85 1.17 1.77 1.17  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.9 -0.085 1.9 0.085 1.665 0.085 1.665 0.49 1.595 0.49 1.595 0.085 1.445 0.085 1.445 0.285 1.31 0.285 1.31 0.085 0.645 0.085 0.645 0.32 0.575 0.32 0.575 0.085 0.33 0.085 0.33 0.21 0.195 0.21 0.195 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 0.7 0.78 0.7 0.78 0.84 0.63 0.84  ;
    END
  END D
  PIN GN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.215 0.42 0.215 0.56 0.06 0.56  ;
    END
  END GN
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.75 0.28 0.75 0.28 0.35 0.045 0.35 0.045 0.215 0.115 0.215 0.115 0.28 0.35 0.28 0.35 0.82 0.115 0.82 0.115 1.065 0.045 1.065  ;
        POLYGON 0.42 0.215 0.49 0.215 0.49 0.945 0.845 0.945 0.845 0.6 0.915 0.6 0.915 1.015 0.42 1.015  ;
        POLYGON 0.96 1.07 0.98 1.07 0.98 0.425 0.95 0.425 0.95 0.29 1.05 0.29 1.05 0.63 1.295 0.63 1.295 0.765 1.05 0.765 1.05 1.205 0.96 1.205  ;
        POLYGON 1.195 0.94 1.365 0.94 1.365 0.47 1.22 0.47 1.22 0.4 1.5 0.4 1.5 1.01 1.195 1.01  ;
  END
END DLL_X2

MACRO FA_X1
  CLASS core ;
  FOREIGN FA_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 3.04 BY 1.4 ;
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.91 0.325 2.985 0.325 2.985 1.065 2.91 1.065  ;
    END
  END S
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.515 0.595 1.515 0.595 1.515 0.665 0.515 0.665  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.25 1.315 0.25 1.175 0.32 1.175 0.32 1.315 0.975 1.315 0.975 1.21 1.11 1.21 1.11 1.315 1.365 1.315 1.365 1.115 1.5 1.115 1.5 1.315 2.315 1.315 2.315 1.025 2.45 1.025 2.45 1.315 2.725 1.315 2.725 0.99 2.795 0.99 2.795 1.315 3.04 1.315 3.04 1.485 0 1.485  ;
    END
  END VDD
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.15 0.13 0.15 0.13 1.25 0.06 1.25  ;
    END
  END CO
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 3.04 -0.085 3.04 0.085 2.795 0.085 2.795 0.445 2.725 0.445 2.725 0.085 2.45 0.085 2.45 0.41 2.315 0.41 2.315 0.085 1.465 0.085 1.465 0.37 1.395 0.37 1.395 0.085 1.075 0.085 1.075 0.23 1.005 0.23 1.005 0.085 0.355 0.085 0.355 0.235 0.22 0.235 0.22 0.085 0 0.085  ;
    END
  END VSS
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.705 0.735 0.925 0.735 0.925 0.765 1.93 0.765 1.93 0.835 0.705 0.835  ;
    END
  END CI
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.33 0.46 1.735 0.46 1.735 0.595 1.65 0.595 1.65 0.7 1.58 0.7 1.58 0.53 0.33 0.53  ;
    END
  END B
  OBS
      LAYER metal1 ;
        POLYGON 0.825 0.15 0.895 0.15 0.895 0.295 1.195 0.295 1.195 0.15 1.265 0.15 1.265 0.365 0.825 0.365  ;
        POLYGON 0.79 1.075 1.3 1.075 1.3 1.15 1.165 1.15 1.165 1.145 0.925 1.145 0.925 1.15 0.79 1.15  ;
        POLYGON 0.265 0.905 1.635 0.905 1.635 1.095 2.12 1.095 2.12 1.25 2.05 1.25 2.05 1.165 1.565 1.165 1.565 0.975 0.695 0.975 0.695 1.185 0.625 1.185 0.625 0.975 0.195 0.975 0.195 0.325 0.625 0.325 0.625 0.15 0.695 0.15 0.695 0.395 0.265 0.395  ;
        POLYGON 2.165 0.365 2.235 0.365 2.235 0.475 2.535 0.475 2.535 0.365 2.605 0.365 2.605 0.545 2.165 0.545  ;
        POLYGON 2.13 0.89 2.64 0.89 2.64 0.965 2.505 0.965 2.505 0.96 2.265 0.96 2.265 0.965 2.13 0.965  ;
        POLYGON 1.975 0.895 1.995 0.895 1.995 0.465 1.975 0.465 1.975 0.33 2.065 0.33 2.065 0.74 2.845 0.74 2.845 0.875 2.775 0.875 2.775 0.81 2.065 0.81 2.065 1.03 1.975 1.03  ;
  END
END FA_X1

MACRO FILLCELL_X1
  CLASS core ;
  FOREIGN FILLCELL_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.19 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.19 1.315 0.19 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.19 -0.085 0.19 0.085 0 0.085  ;
    END
  END VSS
END FILLCELL_X1

MACRO FILLCELL_X16
  CLASS core ;
  FOREIGN FILLCELL_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 3.04 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 3.04 1.315 3.04 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 3.04 -0.085 3.04 0.085 0 0.085  ;
    END
  END VSS
END FILLCELL_X16

MACRO FILLCELL_X2
  CLASS core ;
  FOREIGN FILLCELL_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.38 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.38 1.315 0.38 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.38 -0.085 0.38 0.085 0 0.085  ;
    END
  END VSS
END FILLCELL_X2

MACRO FILLCELL_X32
  CLASS core ;
  FOREIGN FILLCELL_X32 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 6.08 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 6.08 1.315 6.08 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 6.08 -0.085 6.08 0.085 0 0.085  ;
    END
  END VSS
END FILLCELL_X32

MACRO FILLCELL_X4
  CLASS core ;
  FOREIGN FILLCELL_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0 0.085  ;
    END
  END VSS
END FILLCELL_X4

MACRO FILLCELL_X8
  CLASS core ;
  FOREIGN FILLCELL_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.52 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 1.52 1.315 1.52 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.52 -0.085 1.52 0.085 0 0.085  ;
    END
  END VSS
END FILLCELL_X8

MACRO HA_X1
  CLASS core ;
  FOREIGN HA_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.9 BY 1.4 ;
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.615 0.24 0.7 0.24 0.7 0.35 0.825 0.35 0.825 0.96 0.865 0.96 0.865 1.095 0.755 1.095 0.755 0.42 0.615 0.42  ;
    END
  END S
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.19 0.56 0.19 0.7 0.06 0.7  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.42 1.315 0.42 1.02 0.49 1.02 0.49 1.315 1.14 1.315 1.14 1.08 1.21 1.08 1.21 1.315 1.515 1.315 1.515 1.08 1.585 1.08 1.585 1.315 1.9 1.315 1.9 1.485 0 1.485  ;
    END
  END VDD
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.71 1.02 1.77 1.02 1.77 0.285 1.71 0.285 1.71 0.15 1.84 0.15 1.84 1.155 1.71 1.155  ;
    END
  END CO
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.9 -0.085 1.9 0.085 1.59 0.085 1.59 0.27 1.52 0.27 1.52 0.085 1.055 0.085 1.055 0.32 0.985 0.32 0.985 0.085 0.485 0.085 0.485 0.36 0.415 0.36 0.415 0.085 0.11 0.085 0.11 0.36 0.04 0.36 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.905 0.42 1.08 0.42 1.08 0.56 0.905 0.56  ;
    END
  END B
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.765 0.255 0.765 0.255 0.375 0.235 0.375 0.235 0.24 0.325 0.24 0.325 0.485 0.605 0.485 0.605 0.555 0.325 0.555 0.325 0.835 0.115 0.835 0.115 1.095 0.045 1.095  ;
        POLYGON 0.615 1.02 0.685 1.02 0.685 1.16 0.985 1.16 0.985 1.02 1.055 1.02 1.055 1.23 0.615 1.23  ;
        POLYGON 1.145 0.19 1.215 0.19 1.215 0.695 1.705 0.695 1.705 0.765 1.375 0.765 1.375 1.02 1.395 1.02 1.395 1.155 1.305 1.155 1.305 0.765 1.145 0.765  ;
  END
END HA_X1

MACRO INV_X1
  CLASS core ;
  FOREIGN INV_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.38 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.185 0.42 0.185 0.56 0.06 0.56  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.175 0.11 1.175 0.11 1.315 0.38 1.315 0.38 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.38 -0.085 0.38 0.085 0.11 0.085 0.11 0.27 0.04 0.27 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.23 1.115 0.25 1.115 0.25 0.285 0.23 0.285 0.23 0.15 0.32 0.15 0.32 1.25 0.23 1.25  ;
    END
  END ZN
END INV_X1

MACRO INV_X16
  CLASS core ;
  FOREIGN INV_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.615 0.17 0.615 0.17 0.84 0.06 0.84  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.065 0.11 1.065 0.11 1.315 0.385 1.315 0.385 1.24 0.52 1.24 0.52 1.315 0.795 1.315 0.795 1.065 0.865 1.065 0.865 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.865 0.085 0.865 0.48 0.795 0.48 0.795 0.085 0.52 0.085 0.52 0.3 0.385 0.3 0.385 0.085 0.11 0.085 0.11 0.335 0.04 0.335 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.235 0.345 0.305 0.345 0.305 0.685 0.575 0.685 0.575 0.38 0.71 0.38 0.71 0.98 0.575 0.98 0.575 0.845 0.305 0.845 0.305 1.015 0.235 1.015  ;
    END
  END ZN
END INV_X16

MACRO INV_X2
  CLASS core ;
  FOREIGN INV_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.38 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.185 0.42 0.185 0.56 0.06 0.56  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.03 0.11 1.03 0.11 1.315 0.38 1.315 0.38 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.38 -0.085 0.38 0.085 0.11 0.085 0.11 0.195 0.04 0.195 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.23 0.975 0.25 0.975 0.25 0.285 0.23 0.285 0.23 0.15 0.32 0.15 0.32 1.25 0.23 1.25  ;
    END
  END ZN
END INV_X2

MACRO INV_X32
  CLASS core ;
  FOREIGN INV_X32 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.52 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.28 0.185 0.28 0.185 0.655 0.06 0.655  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.055 1.315 0.055 1.065 0.125 1.065 0.125 1.315 0.4 1.315 0.4 1.1 0.535 1.1 0.535 1.315 0.78 1.315 0.78 1.1 0.915 1.1 0.915 1.315 1.16 1.315 1.16 1.1 1.295 1.1 1.295 1.315 1.52 1.315 1.52 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.52 -0.085 1.52 0.085 1.295 0.085 1.295 0.3 1.16 0.3 1.16 0.085 0.915 0.085 0.915 0.3 0.78 0.3 0.78 0.085 0.535 0.085 0.535 0.3 0.4 0.3 0.4 0.085 0.125 0.085 0.125 0.195 0.055 0.195 0.055 0.085 0 0.085  ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.395 0.32 0.395 0.32 0.615 0.62 0.615 0.62 0.395 0.69 0.395 0.69 0.615 1 0.615 1 0.395 1.07 0.395 1.07 0.615 1.38 0.615 1.38 0.395 1.45 0.395 1.45 0.94 1.38 0.94 1.38 0.735 1.105 0.735 1.105 0.94 0.975 0.94 0.975 0.74 0.69 0.74 0.69 0.94 0.62 0.94 0.62 0.74 0.32 0.74 0.32 0.94 0.25 0.94  ;
    END
  END ZN
END INV_X32

MACRO INV_X4
  CLASS core ;
  FOREIGN INV_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.38 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.13 0.42 0.13 0.48 0.19 0.48 0.19 0.615 0.06 0.615  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.065 0.11 1.065 0.11 1.315 0.38 1.315 0.38 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.38 -0.085 0.38 0.085 0.11 0.085 0.11 0.335 0.04 0.335 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.23 0.975 0.255 0.975 0.255 0.425 0.23 0.425 0.23 0.15 0.325 0.15 0.325 1.25 0.23 1.25  ;
    END
  END ZN
END INV_X4

MACRO INV_X8
  CLASS core ;
  FOREIGN INV_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.28 0.185 0.28 0.185 0.605 0.06 0.605  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.055 1.315 0.055 1.065 0.125 1.065 0.125 1.315 0.43 1.315 0.43 1.065 0.5 1.065 0.5 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.5 0.085 0.5 0.335 0.43 0.335 0.43 0.085 0.125 0.085 0.125 0.195 0.055 0.195 0.055 0.085 0 0.085  ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.205 0.32 0.205 0.32 1.015 0.25 1.015  ;
    END
  END ZN
END INV_X8

MACRO LOGIC0_X1
  CLASS core ;
  FOREIGN LOGIC0_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.38 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.195 0.16 0.195 0.16 0.42 0.06 0.42  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.09 1.315 0.09 1.115 0.16 1.115 0.16 1.315 0.38 1.315 0.38 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.38 -0.085 0.38 0.085 0.195 0.085 0.195 0.11 0.06 0.11 0.06 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.075 0.69 0.31 0.69 0.31 0.76 0.21 0.76 0.21 1.03 0.075 1.03  ;
  END
END LOGIC0_X1

MACRO LOGIC1_X1
  CLASS core ;
  FOREIGN LOGIC1_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.38 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.175 0.56 0.175 1.19 0.06 1.19  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.15 1.315 0.15 1.255 0.22 1.255 0.22 1.315 0.38 1.315 0.38 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.38 -0.085 0.38 0.085 0.195 0.085 0.195 0.145 0.125 0.145 0.125 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.11 0.23 0.335 0.23 0.335 0.44 0.22 0.44 0.22 0.3 0.11 0.3  ;
  END
END LOGIC1_X1

MACRO MUX2_X1
  CLASS core ;
  FOREIGN MUX2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.33 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.2 0.165 1.27 0.165 1.27 1.195 1.2 1.195  ;
    END
  END Z
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.17 0.42 0.32 0.42 0.32 0.56 0.17 0.56  ;
    END
  END S
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.59 0.29 0.7 0.29 0.7 0.805 1 0.805 1 0.875 0.59 0.875  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.24 1.315 0.24 1.075 0.31 1.075 0.31 1.315 1.005 1.315 1.005 1.12 1.075 1.12 1.075 1.315 1.33 1.315 1.33 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.33 -0.085 1.33 0.085 1.075 0.085 1.075 0.285 1.005 0.285 1.005 0.085 0.31 0.085 0.31 0.195 0.24 0.195 0.24 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.765 0.42 0.89 0.42 0.89 0.7 0.765 0.7  ;
    END
  END B
  OBS
      LAYER metal1 ;
        POLYGON 0.105 0.88 0.39 0.88 0.39 0.95 0.125 0.95 0.125 1.105 0.035 1.105 0.035 0.165 0.125 0.165 0.125 0.3 0.105 0.3  ;
        POLYGON 0.44 1.075 0.51 1.075 0.51 1.18 0.81 1.18 0.81 1.075 0.88 1.075 0.88 1.25 0.44 1.25  ;
        POLYGON 0.525 0.94 1.065 0.94 1.065 0.875 1.135 0.875 1.135 1.01 0.725 1.01 0.725 1.115 0.59 1.115 0.59 1.01 0.455 1.01 0.455 0.155 0.73 0.155 0.73 0.225 0.525 0.225  ;
  END
END MUX2_X1

MACRO MUX2_X2
  CLASS core ;
  FOREIGN MUX2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.33 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.2 0.165 1.275 0.165 1.275 1.145 1.2 1.145  ;
    END
  END Z
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.17 0.42 0.32 0.42 0.32 0.56 0.17 0.56  ;
    END
  END S
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.59 0.29 0.7 0.29 0.7 0.845 1 0.845 1 0.915 0.59 0.915  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.24 1.315 0.24 1.08 0.31 1.08 0.31 1.315 1.015 1.315 1.015 1.115 1.085 1.115 1.085 1.315 1.33 1.315 1.33 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.33 -0.085 1.33 0.085 1.075 0.085 1.075 0.195 1.005 0.195 1.005 0.085 0.31 0.085 0.31 0.195 0.24 0.195 0.24 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.765 0.42 0.89 0.42 0.89 0.7 0.765 0.7  ;
    END
  END B
  OBS
      LAYER metal1 ;
        POLYGON 0.105 0.885 0.39 0.885 0.39 0.955 0.125 0.955 0.125 1.11 0.035 1.11 0.035 0.165 0.125 0.165 0.125 0.3 0.105 0.3  ;
        POLYGON 0.4 1.115 0.535 1.115 0.535 1.145 0.93 1.145 0.93 1.215 0.4 1.215  ;
        POLYGON 0.525 0.98 1.065 0.98 1.065 0.885 1.135 0.885 1.135 1.05 0.725 1.05 0.725 1.08 0.59 1.08 0.59 1.05 0.455 1.05 0.455 0.155 0.73 0.155 0.73 0.225 0.525 0.225  ;
  END
END MUX2_X2

MACRO NAND2_X1
  CLASS core ;
  FOREIGN NAND2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.175 0.11 1.175 0.11 1.315 0.415 1.315 0.415 1.175 0.485 1.175 0.485 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.28 0.355 0.28 0.355 0.42 0.25 0.42  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.11 0.085 0.11 0.23 0.04 0.23 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.185 0.42 0.185 0.56 0.06 0.56  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.235 0.98 0.42 0.98 0.42 0.15 0.49 0.15 0.49 1.05 0.32 1.05 0.32 1.25 0.235 1.25  ;
    END
  END ZN
END NAND2_X1

MACRO NAND2_X2
  CLASS core ;
  FOREIGN NAND2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.03 0.11 1.03 0.11 1.315 0.415 1.315 0.415 1.03 0.485 1.03 0.485 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.28 0.355 0.28 0.355 0.505 0.25 0.505  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.11 0.085 0.11 0.195 0.04 0.195 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.28 0.185 0.28 0.185 0.505 0.06 0.505  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.235 0.895 0.42 0.895 0.42 0.245 0.51 0.245 0.51 0.965 0.305 0.965 0.305 1.25 0.235 1.25  ;
    END
  END ZN
END NAND2_X2

MACRO NAND2_X4
  CLASS core ;
  FOREIGN NAND2_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.08 1.315 0.08 1.03 0.15 1.03 0.15 1.315 0.455 1.315 0.455 1.17 0.525 1.17 0.525 1.315 0.835 1.315 0.835 1.03 0.905 1.03 0.905 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.535 0.875 0.735 0.875 0.735 0.945 0.535 0.945  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.91 0.085 0.91 0.375 0.84 0.375 0.84 0.085 0.15 0.085 0.15 0.375 0.08 0.375 0.08 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.19 0.43 0.25 0.43 0.25 0.15 0.775 0.15 0.775 0.545 0.705 0.545 0.705 0.22 0.32 0.22 0.32 0.565 0.19 0.565  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.345 1.01 0.75 1.01 0.75 1.08 0.345 1.08 0.345 1.25 0.275 1.25 0.275 0.74 0.42 0.74 0.42 0.285 0.525 0.285 0.525 0.81 0.345 0.81  ;
    END
  END ZN
END NAND2_X4

MACRO NAND3_X1
  CLASS core ;
  FOREIGN NAND3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.175 0.11 1.175 0.11 1.315 0.42 1.315 0.42 1.175 0.49 1.175 0.49 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.28 0.13 0.28 0.13 0.475 0.215 0.475 0.215 0.61 0.06 0.61  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.28 0.545 0.28 0.545 0.42 0.44 0.42  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.11 0.085 0.11 0.195 0.04 0.195 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.28 0.375 0.28 0.375 0.42 0.25 0.42  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.235 0.98 0.61 0.98 0.61 0.155 0.68 0.155 0.68 1.25 0.61 1.25 0.61 1.05 0.32 1.05 0.32 1.25 0.235 1.25  ;
    END
  END ZN
END NAND3_X1

MACRO NAND3_X2
  CLASS core ;
  FOREIGN NAND3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.065 0.11 1.065 0.11 1.315 0.385 1.315 0.385 1.24 0.52 1.24 0.52 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.28 0.19 0.28 0.19 0.59 0.06 0.59  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.28 0.545 0.28 0.545 0.59 0.44 0.59  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.11 0.085 0.11 0.195 0.04 0.195 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.84 0.415 0.84 0.415 0.98 0.25 0.98  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2 1.075 0.61 1.075 0.61 0.185 0.7 0.185 0.7 1.145 0.2 1.145  ;
    END
  END ZN
END NAND3_X2

MACRO NAND3_X4
  CLASS core ;
  FOREIGN NAND3_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.33 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.065 0.11 1.065 0.11 1.315 0.385 1.315 0.385 1.24 0.52 1.24 0.52 1.315 0.77 1.315 0.77 1.24 0.905 1.24 0.905 1.315 1.18 1.315 1.18 0.74 1.25 0.74 1.25 1.315 1.33 1.315 1.33 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.15 0.545 0.175 0.545 0.175 0.15 1.09 0.15 1.09 0.575 1.18 0.575 1.18 0.645 1.02 0.645 1.02 0.42 1.01 0.42 1.01 0.22 0.245 0.22 0.245 0.68 0.15 0.68  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.74 0.615 0.81 0.615 0.81 0.84 0.89 0.84 0.89 0.98 0.74 0.98  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.33 -0.085 1.33 0.085 1.25 0.085 1.25 0.43 1.18 0.43 1.18 0.085 0.11 0.085 0.11 0.43 0.04 0.43 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.31 0.575 0.44 0.575 0.44 0.285 0.945 0.285 0.945 0.545 0.955 0.545 0.955 0.68 0.875 0.68 0.875 0.355 0.51 0.355 0.51 0.645 0.31 0.645  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2 0.915 0.335 0.915 0.335 1.045 0.605 1.045 0.605 0.42 0.675 0.42 0.675 1.045 0.96 1.045 0.96 0.91 1.095 0.91 1.095 1.12 0.2 1.12  ;
    END
  END ZN
END NAND3_X4

MACRO NAND4_X1
  CLASS core ;
  FOREIGN NAND4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.175 0.11 1.175 0.11 1.315 0.42 1.315 0.42 1.175 0.49 1.175 0.49 1.315 0.795 1.315 0.795 1.175 0.865 1.175 0.865 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.28 0.375 0.28 0.375 0.46 0.25 0.46  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 0.28 0.735 0.28 0.735 0.46 0.63 0.46  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.11 0.085 0.11 0.195 0.04 0.195 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.28 0.565 0.28 0.565 0.46 0.44 0.46  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.28 0.185 0.28 0.185 0.46 0.06 0.46  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.235 0.98 0.8 0.98 0.8 0.2 0.87 0.2 0.87 1.05 0.675 1.05 0.675 1.25 0.605 1.25 0.605 1.05 0.32 1.05 0.32 1.25 0.235 1.25  ;
    END
  END ZN
END NAND4_X1

MACRO NAND4_X2
  CLASS core ;
  FOREIGN NAND4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.065 0.11 1.065 0.11 1.315 0.385 1.315 0.385 1.24 0.52 1.24 0.52 1.315 0.795 1.315 0.795 1.205 0.865 1.205 0.865 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.28 0.32 0.28 0.32 0.545 0.405 0.545 0.405 0.68 0.25 0.68  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 0.84 0.76 0.84 0.76 0.98 0.63 0.98  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.11 0.085 0.11 0.195 0.04 0.195 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.28 0.595 0.28 0.595 0.68 0.525 0.68 0.525 0.42 0.44 0.42  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.28 0.13 0.28 0.13 0.705 0.19 0.705 0.19 0.84 0.06 0.84  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2 1.045 0.825 1.045 0.825 0.555 0.8 0.555 0.8 0.275 0.895 0.275 0.895 1.115 0.2 1.115  ;
    END
  END ZN
END NAND4_X2

MACRO NAND4_X4
  CLASS core ;
  FOREIGN NAND4_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.71 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.08 1.315 0.08 1.205 0.15 1.205 0.15 1.315 0.455 1.315 0.455 1.205 0.525 1.205 0.525 1.315 0.835 1.315 0.835 1.205 0.905 1.205 0.905 1.315 1.215 1.315 1.215 1.205 1.285 1.205 1.285 1.315 1.595 1.315 1.595 1.065 1.665 1.065 1.665 1.315 1.71 1.315 1.71 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.345 0.56 1.405 0.56 1.405 0.7 1.2 0.7 1.2 0.635 0.48 0.635 0.48 0.645 0.345 0.645  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.725 0.7 0.89 0.7 0.89 0.84 0.725 0.84  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.71 -0.085 1.71 0.085 1.665 0.085 1.665 0.195 1.595 0.195 1.595 0.085 0.15 0.085 0.15 0.195 0.08 0.195 0.08 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.84 0.635 0.84 0.635 0.91 1.24 0.91 1.24 0.98 0.44 0.98  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.195 0.41 1.39 0.41 1.39 0.28 1.56 0.28 1.56 0.68 1.49 0.68 1.49 0.48 0.265 0.48 0.265 0.68 0.195 0.68  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.13 1.045 1.51 1.045 1.51 1.115 0.06 1.115 0.06 0.27 0.94 0.27 0.94 0.34 0.13 0.34  ;
    END
  END ZN
END NAND4_X4

MACRO NOR2_X1
  CLASS core ;
  FOREIGN NOR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.205 0.11 1.205 0.11 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.96 0.355 0.96 0.355 1.12 0.25 1.12  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.505 0.085 0.505 0.215 0.435 0.215 0.435 0.085 0.11 0.085 0.11 0.27 0.04 0.27 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.96 0.185 0.96 0.185 1.12 0.06 1.12  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.235 0.15 0.305 0.15 0.305 0.28 0.51 0.28 0.51 1.22 0.42 1.22 0.42 0.35 0.235 0.35  ;
    END
  END ZN
END NOR2_X1

MACRO NOR2_X2
  CLASS core ;
  FOREIGN NOR2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.055 1.315 0.055 1.065 0.125 1.065 0.125 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.385 0.28 0.51 0.28 0.51 0.425 0.385 0.425  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.5 0.085 0.5 0.195 0.43 0.195 0.43 0.085 0.125 0.085 0.125 0.195 0.055 0.195 0.055 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.28 0.185 0.28 0.185 0.425 0.06 0.425  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.165 0.32 0.165 0.32 0.49 0.5 0.49 0.5 1.165 0.43 1.165 0.43 0.56 0.25 0.56  ;
    END
  END ZN
END NOR2_X2

MACRO NOR2_X4
  CLASS core ;
  FOREIGN NOR2_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.02 0.11 1.02 0.11 1.315 0.795 1.315 0.795 1.02 0.865 1.02 0.865 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.49 0.28 0.7 0.28 0.7 0.42 0.56 0.42 0.56 0.775 0.49 0.775  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.505 0.085 0.505 0.195 0.435 0.195 0.435 0.085 0.13 0.085 0.13 0.335 0.06 0.335 0.06 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.15 0.715 0.245 0.715 0.245 1.18 0.63 1.18 0.63 0.715 0.76 0.715 0.76 0.85 0.7 0.85 0.7 1.25 0.175 1.25 0.175 0.85 0.15 0.85  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.205 0.32 0.205 0.32 0.41 0.42 0.41 0.42 0.875 0.52 0.875 0.52 1.085 0.35 1.085 0.35 0.48 0.25 0.48  ;
    END
  END ZN
END NOR2_X4

MACRO NOR3_X1
  CLASS core ;
  FOREIGN NOR3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.02 0.11 1.02 0.11 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.19 0.56 0.19 0.7 0.06 0.7  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.85 0.545 0.85 0.545 1.12 0.44 1.12  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.49 0.085 0.49 0.27 0.42 0.27 0.42 0.085 0.11 0.085 0.11 0.27 0.04 0.27 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.85 0.375 0.85 0.375 1.12 0.25 1.12  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.235 0.15 0.32 0.15 0.32 0.35 0.61 0.35 0.61 0.15 0.68 0.15 0.68 1.25 0.61 1.25 0.61 0.42 0.235 0.42  ;
    END
  END ZN
END NOR3_X1

MACRO NOR3_X2
  CLASS core ;
  FOREIGN NOR3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.065 0.11 1.065 0.11 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.63 0.185 0.63 0.185 0.84 0.06 0.84  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.58 0.56 0.58 0.56 0.715 0.51 0.715 0.51 0.84 0.44 0.84  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.485 0.085 0.485 0.195 0.415 0.195 0.415 0.085 0.11 0.085 0.11 0.195 0.04 0.195 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.63 0.375 0.63 0.375 0.84 0.25 0.84  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.61 0.76 0.63 0.76 0.63 0.33 0.235 0.33 0.235 0.165 0.305 0.165 0.305 0.26 0.61 0.26 0.61 0.165 0.7 0.165 0.7 1.035 0.61 1.035  ;
    END
  END ZN
END NOR3_X2

MACRO NOR3_X4
  CLASS core ;
  FOREIGN NOR3_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.33 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.205 0.11 1.205 0.11 1.315 1.175 1.315 1.175 1.205 1.245 1.205 1.245 1.315 1.33 1.315 1.33 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.15 0.63 0.245 0.63 0.245 1.09 1.01 1.09 1.01 0.84 1.05 0.84 1.05 0.63 1.14 0.63 1.14 0.765 1.12 0.765 1.12 1.16 0.175 1.16 0.175 0.765 0.15 0.765  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.71 0.42 0.89 0.42 0.89 0.56 0.78 0.56 0.78 0.61 0.71 0.61  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.33 -0.085 1.33 0.085 0.525 0.085 0.525 0.16 0.39 0.16 0.39 0.085 0.11 0.085 0.11 0.335 0.04 0.335 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.34 0.63 0.41 0.63 0.41 0.955 0.82 0.955 0.82 0.665 0.985 0.665 0.985 0.735 0.89 0.735 0.89 1.025 0.34 1.025  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.645 0.7 0.71 0.7 0.71 0.86 0.575 0.86 0.575 0.35 0.2 0.35 0.2 0.28 0.71 0.28 0.71 0.35 0.645 0.35  ;
    END
  END ZN
END NOR3_X4

MACRO NOR4_X1
  CLASS core ;
  FOREIGN NOR4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.065 0.11 1.065 0.11 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.83 0.375 0.83 0.375 0.98 0.25 0.98  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 0.83 0.735 0.83 0.735 0.98 0.63 0.98  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.865 0.085 0.865 0.27 0.795 0.27 0.795 0.085 0.49 0.085 0.49 0.27 0.42 0.27 0.42 0.085 0.11 0.085 0.11 0.27 0.04 0.27 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.83 0.565 0.83 0.565 0.98 0.44 0.98  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.19 0.56 0.19 0.7 0.06 0.7  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.235 0.15 0.32 0.15 0.32 0.35 0.605 0.35 0.605 0.15 0.675 0.15 0.675 0.35 0.87 0.35 0.87 1.23 0.8 1.23 0.8 0.42 0.235 0.42  ;
    END
  END ZN
END NOR4_X1

MACRO NOR4_X2
  CLASS core ;
  FOREIGN NOR4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.065 0.11 1.065 0.11 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.42 0.375 0.42 0.375 0.56 0.25 0.56  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 0.505 0.74 0.505 0.74 0.7 0.63 0.7  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.865 0.085 0.865 0.195 0.795 0.195 0.795 0.085 0.49 0.085 0.49 0.195 0.42 0.195 0.42 0.085 0.11 0.085 0.11 0.195 0.04 0.195 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.505 0.565 0.505 0.565 0.7 0.44 0.7  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.185 0.42 0.185 0.56 0.06 0.56  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.8 0.725 0.805 0.725 0.805 0.42 0.44 0.42 0.44 0.35 0.235 0.35 0.235 0.165 0.305 0.165 0.305 0.28 0.605 0.28 0.605 0.165 0.675 0.165 0.675 0.35 0.875 0.35 0.875 1 0.8 1  ;
    END
  END ZN
END NOR4_X2

MACRO NOR4_X4
  CLASS core ;
  FOREIGN NOR4_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.71 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.08 1.315 0.08 1.065 0.15 1.065 0.15 1.315 1.6 1.315 1.6 1.065 1.67 1.065 1.67 1.315 1.71 1.315 1.71 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.38 0.505 0.45 0.505 0.45 1.015 1.295 1.015 1.295 0.505 1.365 0.505 1.365 1.085 0.38 1.085  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.81 0.42 0.89 0.42 0.89 0.56 0.81 0.56  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.71 -0.085 1.71 0.085 1.665 0.085 1.665 0.195 1.595 0.195 1.595 0.085 1.32 0.085 1.32 0.16 1.185 0.16 1.185 0.085 0.94 0.085 0.94 0.16 0.805 0.16 0.805 0.085 0.56 0.085 0.56 0.16 0.425 0.16 0.425 0.085 0.185 0.085 0.185 0.16 0.05 0.16 0.05 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.57 0.505 0.64 0.505 0.64 0.875 1.11 0.875 1.11 0.505 1.18 0.505 1.18 0.945 0.57 0.945  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.19 0.505 0.285 0.505 0.285 1.155 1.465 1.155 1.465 0.505 1.56 0.505 1.56 0.64 1.535 0.64 1.535 1.225 0.215 1.225 0.215 0.64 0.19 0.64  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.81 0.665 0.97 0.665 0.97 0.35 0.13 0.35 0.13 0.42 0.055 0.42 0.055 0.265 0.265 0.265 0.265 0.165 0.335 0.165 0.335 0.265 0.645 0.265 0.645 0.165 0.715 0.165 0.715 0.265 1.025 0.265 1.025 0.165 1.095 0.165 1.095 0.265 1.405 0.265 1.405 0.165 1.475 0.165 1.475 0.35 1.04 0.35 1.04 0.735 0.81 0.735  ;
    END
  END ZN
END NOR4_X4

MACRO OAI211_X1
  CLASS core ;
  FOREIGN OAI211_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.575 0.41 0.63 0.41 0.63 0.28 0.7 0.28 0.7 0.545 0.575 0.545  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.08 1.315 0.08 1.175 0.15 1.175 0.15 1.315 0.645 1.315 0.645 1.175 0.715 1.175 0.715 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.905 0.085 0.905 0.325 0.835 0.325 0.835 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.765 0.42 0.89 0.42 0.89 0.56 0.765 0.56  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.285 0.335 0.285 0.335 1.04 0.905 1.04 0.905 1.25 0.835 1.25 0.835 1.11 0.53 1.11 0.53 1.25 0.46 1.25 0.46 1.11 0.25 1.11  ;
    END
  END ZN
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.185 0.42 0.185 0.56 0.06 0.56  ;
    END
  END C2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4 0.42 0.51 0.42 0.51 0.56 0.4 0.56  ;
    END
  END C1
  OBS
      LAYER metal1 ;
        POLYGON 0.085 0.15 0.525 0.15 0.525 0.325 0.455 0.325 0.455 0.22 0.155 0.22 0.155 0.325 0.085 0.325  ;
  END
END OAI211_X1

MACRO OAI211_X2
  CLASS core ;
  FOREIGN OAI211_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.575 0.455 0.63 0.455 0.63 0.42 0.7 0.42 0.7 0.59 0.575 0.59  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.07 1.315 0.07 1.005 0.14 1.005 0.14 1.315 0.635 1.315 0.635 1.005 0.705 1.005 0.705 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.895 0.085 0.895 0.195 0.825 0.195 0.825 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.765 0.28 0.89 0.28 0.89 0.59 0.765 0.59  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.325 0.325 0.325 0.325 0.87 0.895 0.87 0.895 1.225 0.825 1.225 0.825 0.94 0.515 0.94 0.515 1.225 0.445 1.225 0.445 0.94 0.25 0.94  ;
    END
  END ZN
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.185 0.42 0.185 0.59 0.06 0.59  ;
    END
  END C2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.39 0.56 0.51 0.56 0.51 0.7 0.39 0.7  ;
    END
  END C1
  OBS
      LAYER metal1 ;
        POLYGON 0.04 0.15 0.515 0.15 0.515 0.425 0.445 0.425 0.445 0.22 0.04 0.22  ;
  END
END OAI211_X2

MACRO OAI211_X4
  CLASS core ;
  FOREIGN OAI211_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.71 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.965 0.395 1.56 0.395 1.56 0.59 1.49 0.59 1.49 0.465 1.08 0.465 1.08 0.59 0.965 0.59  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.05 1.315 0.05 1.065 0.12 1.065 0.12 1.315 0.815 1.315 0.815 1.205 0.885 1.205 0.885 1.315 1.19 1.315 1.19 1.065 1.26 1.065 1.26 1.315 1.71 1.315 1.71 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.71 -0.085 1.71 0.085 1.26 0.085 1.26 0.195 1.19 0.195 1.19 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.145 0.53 1.27 0.53 1.27 0.7 1.145 0.7  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4 1.05 0.795 1.05 0.795 0.465 0.21 0.465 0.21 0.36 0.725 0.36 0.725 0.395 0.865 0.395 0.865 0.975 1.07 0.975 1.07 1.25 1 1.25 1 1.12 0.4 1.12  ;
    END
  END ZN
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1 0.56 0.73 0.56 0.73 0.7 0.63 0.7 0.63 0.63 0.1 0.63  ;
    END
  END C2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.7 0.39 0.7 0.39 0.84 0.25 0.84  ;
    END
  END C1
  OBS
      LAYER metal1 ;
        POLYGON 0.055 0.15 0.875 0.15 0.875 0.26 1.675 0.26 1.675 0.33 0.805 0.33 0.805 0.22 0.125 0.22 0.125 0.425 0.055 0.425  ;
  END
END OAI211_X4

MACRO OAI21_X1
  CLASS core ;
  FOREIGN OAI21_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.575 0.7 0.7 0.7 0.7 0.84 0.575 0.84  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.065 1.315 0.065 1.205 0.135 1.205 0.135 1.315 0.63 1.315 0.63 1.145 0.7 1.145 0.7 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.385 0.56 0.51 0.56 0.51 0.7 0.385 0.7  ;
    END
  END B1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.7 0.085 0.7 0.365 0.63 0.365 0.63 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.185 0.56 0.185 0.7 0.06 0.7  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.285 0.32 0.285 0.32 1.085 0.51 1.085 0.51 1.22 0.25 1.22  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.07 0.15 0.51 0.15 0.51 0.365 0.44 0.365 0.44 0.22 0.14 0.22 0.14 0.365 0.07 0.365  ;
  END
END OAI21_X1

MACRO OAI21_X2
  CLASS core ;
  FOREIGN OAI21_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.575 0.42 0.7 0.42 0.7 0.56 0.575 0.56  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.065 1.315 0.065 1.03 0.135 1.03 0.135 1.315 0.63 1.315 0.63 1.03 0.7 1.03 0.7 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.385 0.42 0.51 0.42 0.51 0.56 0.385 0.56  ;
    END
  END B1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.7 0.085 0.7 0.235 0.63 0.235 0.63 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.185 0.42 0.185 0.56 0.06 0.56  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.285 0.32 0.285 0.32 0.975 0.51 0.975 0.51 1.25 0.44 1.25 0.44 1.045 0.25 1.045  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.035 0.15 0.545 0.15 0.545 0.22 0.035 0.22  ;
  END
END OAI21_X2

MACRO OAI21_X4
  CLASS core ;
  FOREIGN OAI21_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.33 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.82 0.84 0.93 0.84 0.93 0.58 1 0.58 1 0.98 0.82 0.98  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.44 1.315 0.44 1.205 0.51 1.205 0.51 1.315 1.01 1.315 1.01 1.065 1.08 1.065 1.08 1.315 1.33 1.315 1.33 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2 0.56 0.32 0.56 0.32 0.625 0.845 0.625 0.845 0.695 0.32 0.695 0.32 0.7 0.2 0.7  ;
    END
  END B1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.33 -0.085 1.33 0.085 1.08 0.085 1.08 0.38 1.01 0.38 1.01 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.84 0.36 0.84 0.36 0.76 0.43 0.76 0.43 0.98 0.25 0.98  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.135 1.045 0.925 1.045 0.925 1.115 0.06 1.115 0.06 0.325 0.735 0.325 0.735 0.395 0.135 0.395  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.035 0.15 0.89 0.15 0.89 0.445 1.2 0.445 1.2 0.15 1.27 0.15 1.27 0.515 0.82 0.515 0.82 0.22 0.035 0.22  ;
  END
END OAI21_X4

MACRO OAI221_X1
  CLASS core ;
  FOREIGN OAI221_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.55 0.42 0.7 0.42 0.7 0.56 0.55 0.56  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.175 0.11 1.175 0.11 1.315 0.605 1.315 0.605 1.175 0.675 1.175 0.675 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.93 0.375 0.93 0.375 1.065 0.32 1.065 0.32 1.12 0.25 1.12  ;
    END
  END B1
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.425 1.115 0.44 1.115 0.44 0.98 0.805 0.98 0.805 0.285 0.875 0.285 0.875 0.99 1.055 0.99 1.055 1.19 0.985 1.19 0.985 1.06 0.51 1.06 0.51 1.25 0.425 1.25  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.94 0.7 1.08 0.7 1.08 0.84 0.94 0.84  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.295 0.085 0.295 0.325 0.225 0.325 0.225 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.215 0.56 0.215 0.7 0.06 0.7  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 0.7 0.74 0.7 0.74 0.84 0.63 0.84  ;
    END
  END C2
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.285 0.115 0.285 0.115 0.39 0.415 0.39 0.415 0.285 0.485 0.285 0.485 0.46 0.045 0.46  ;
        POLYGON 0.615 0.15 1.055 0.15 1.055 0.325 0.985 0.325 0.985 0.22 0.685 0.22 0.685 0.325 0.615 0.325  ;
  END
END OAI221_X1

MACRO OAI221_X2
  CLASS core ;
  FOREIGN OAI221_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.42 0.565 0.42 0.565 0.59 0.44 0.59  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.065 0.11 1.065 0.11 1.315 0.605 1.315 0.605 1.205 0.675 1.205 0.675 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.76 0.38 0.76 0.38 0.895 0.32 0.895 0.32 0.98 0.25 0.98  ;
    END
  END B1
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.39 1.045 0.81 1.045 0.81 0.325 0.88 0.325 0.88 0.98 1.06 0.98 1.06 1.12 0.39 1.12  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.945 0.7 1.08 0.7 1.08 0.84 0.945 0.84  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.295 0.085 0.295 0.195 0.225 0.195 0.225 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.25 0.42 0.25 0.56 0.06 0.56  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 0.42 0.745 0.42 0.745 0.59 0.63 0.59  ;
    END
  END C2
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.15 0.115 0.15 0.115 0.26 0.52 0.26 0.52 0.33 0.045 0.33  ;
        POLYGON 0.585 0.165 1.06 0.165 1.06 0.44 0.99 0.44 0.99 0.235 0.585 0.235  ;
  END
END OAI221_X2

MACRO OAI221_X4
  CLASS core ;
  FOREIGN OAI221_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.28 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.135 0.49 1.27 0.49 1.27 0.7 1.135 0.7  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.495 1.315 0.495 1.065 0.565 1.065 0.565 1.315 1.27 1.315 1.27 1.065 1.34 1.065 1.34 1.315 2.03 1.315 2.03 1.065 2.1 1.065 2.1 1.315 2.28 1.315 2.28 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.7 0.69 1.84 0.69 1.84 0.84 1.7 0.84  ;
    END
  END B1
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.105 0.925 1.755 0.925 1.755 0.995 0.035 0.995 0.035 0.15 0.13 0.15 0.13 0.35 0.915 0.35 0.915 0.42 0.105 0.42  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.17 0.565 0.7 0.565 0.7 0.705 0.8 0.705 0.8 0.84 0.63 0.84 0.63 0.635 0.17 0.635  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.28 -0.085 2.28 0.085 1.99 0.085 1.99 0.195 1.92 0.195 1.92 0.085 1.615 0.085 1.615 0.195 1.545 0.195 1.545 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.405 0.555 2.03 0.555 2.03 0.84 1.96 0.84 1.96 0.625 1.54 0.625 1.54 0.69 1.405 0.69  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.7 0.42 0.7 0.42 0.84 0.25 0.84  ;
    END
  END C2
  OBS
      LAYER metal1 ;
        POLYGON 0.215 0.15 1.265 0.15 1.265 0.22 0.215 0.22  ;
        POLYGON 0.98 0.285 2.18 0.285 2.18 0.425 0.98 0.425  ;
  END
END OAI221_X4

MACRO OAI222_X1
  CLASS core ;
  FOREIGN OAI222_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.52 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.31 1.315 0.31 1.1 0.38 1.1 0.38 1.315 1.38 1.315 1.38 0.845 1.45 0.845 1.45 1.315 1.52 1.315 1.52 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.8 0.7 0.89 0.7 0.89 0.84 0.8 0.84  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.01 0.56 1.08 0.56 1.08 0.7 1.01 0.7  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.28 0.42 1.46 0.42 1.46 0.565 1.28 0.565  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.695 1.1 0.765 1.1 0.765 1.18 1.01 1.18 1.01 0.765 1.145 0.765 1.145 0.42 1.1 0.42 1.1 0.285 1.215 0.285 1.215 0.835 1.08 0.835 1.08 1.25 0.695 1.25  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.595 0.735 0.735 0.735 0.735 0.87 0.595 0.87  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.52 -0.085 1.52 0.085 0.59 0.085 0.59 0.325 0.52 0.325 0.52 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.7 0.295 0.7 0.295 0.84 0.06 0.84  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.42 0.7 0.51 0.7 0.51 0.84 0.42 0.84  ;
    END
  END C2
  OBS
      LAYER metal1 ;
        POLYGON 0.34 0.285 0.41 0.285 0.41 0.39 0.71 0.39 0.71 0.285 0.78 0.285 0.78 0.46 0.34 0.46  ;
        POLYGON 0.125 0.965 0.945 0.965 0.945 1.115 0.875 1.115 0.875 1.035 0.195 1.035 0.195 1.115 0.125 1.115  ;
        POLYGON 0.15 0.285 0.22 0.285 0.22 0.525 0.875 0.525 0.875 0.15 1.35 0.15 1.35 0.325 1.28 0.325 1.28 0.22 0.97 0.22 0.97 0.325 0.945 0.325 0.945 0.595 0.15 0.595  ;
  END
END OAI222_X1

MACRO OAI222_X2
  CLASS core ;
  FOREIGN OAI222_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.52 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.27 1.315 0.27 1.065 0.34 1.065 0.34 1.315 1.38 1.315 1.38 1.065 1.45 1.065 1.45 1.315 1.52 1.315 1.52 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.765 0.56 0.89 0.56 0.89 0.7 0.765 0.7  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.98 0.56 1.08 0.56 1.08 0.75 0.98 0.75  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.28 0.42 1.46 0.42 1.46 0.59 1.28 0.59  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.625 1.095 1.145 1.095 1.145 0.43 1.03 0.43 1.03 0.36 1.215 0.36 1.215 0.98 1.27 0.98 1.27 1.165 0.625 1.165  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.575 0.7 0.7 0.7 0.7 0.84 0.575 0.84  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.52 -0.085 1.52 0.085 0.59 0.085 0.59 0.16 0.455 0.16 0.455 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.26 0.56 0.26 0.7 0.06 0.7  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.385 0.56 0.51 0.56 0.51 0.7 0.385 0.7  ;
    END
  END C2
  OBS
      LAYER metal1 ;
        POLYGON 0.27 0.36 0.78 0.36 0.78 0.43 0.27 0.43  ;
        POLYGON 0.09 0.93 0.945 0.93 0.945 1 0.16 1 0.16 1.205 0.09 1.205  ;
        POLYGON 0.08 0.225 1.35 0.225 1.35 0.295 0.08 0.295  ;
  END
END OAI222_X2

MACRO OAI222_X4
  CLASS core ;
  FOREIGN OAI222_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.66 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.065 0.11 1.065 0.11 1.315 0.795 1.315 0.795 1.205 0.865 1.205 0.865 1.315 1.555 1.315 1.555 1.205 1.625 1.205 1.625 1.315 2.12 1.315 2.12 1.205 2.19 1.205 2.19 1.315 2.66 1.315 2.66 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.01 0.76 1.165 0.76 1.165 0.895 1.08 0.895 1.08 0.98 1.01 0.98  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.86 0.625 2.465 0.625 2.465 0.98 2.34 0.98 2.34 0.695 1.86 0.695  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.96 0.76 2.11 0.76 2.11 0.895 2.03 0.895 2.03 0.98 1.96 0.98  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.795 1.05 2.605 1.05 2.605 1.12 0.39 1.12 0.39 1.05 1.2 1.05 1.2 0.98 1.725 0.98 1.725 0.285 1.815 0.285 1.815 0.355 2.5 0.355 2.5 0.15 2.57 0.15 2.57 0.425 1.795 0.425  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.56 0.32 0.56 0.32 0.63 0.44 0.63 0.44 0.7 0.25 0.7  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.66 -0.085 2.66 0.085 0.68 0.085 0.68 0.195 0.61 0.195 0.61 0.085 0.3 0.085 0.3 0.195 0.23 0.195 0.23 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.885 0.56 1.65 0.56 1.65 0.7 1.48 0.7 1.48 0.63 0.885 0.63  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.115 0.42 0.51 0.42 0.51 0.49 0.82 0.49 0.82 0.56 0.44 0.56 0.44 0.49 0.185 0.49 0.185 0.59 0.115 0.59  ;
    END
  END C2
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.15 0.115 0.15 0.115 0.285 1.66 0.285 1.66 0.355 0.045 0.355  ;
        POLYGON 0.96 0.15 2.415 0.15 2.415 0.22 0.96 0.22  ;
  END
END OAI222_X4

MACRO OAI22_X1
  CLASS core ;
  FOREIGN OAI22_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.205 0.11 1.205 0.11 1.315 0.795 1.315 0.795 1.205 0.865 1.205 0.865 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.7 0.35 0.7 0.35 0.84 0.25 0.84  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.405 0.595 0.6 0.595 0.6 0.665 0.405 0.665  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.295 0.085 0.295 0.365 0.225 0.365 0.225 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.7 0.185 0.7 0.185 0.84 0.06 0.84  ;
    END
  END B2
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 0.96 0.785 0.96 0.785 1.12 0.63 1.12  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.425 0.825 0.665 0.825 0.665 0.42 0.615 0.42 0.615 0.285 0.735 0.285 0.735 0.895 0.51 0.895 0.51 1.22 0.425 1.22  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.285 0.115 0.285 0.115 0.43 0.425 0.43 0.425 0.15 0.87 0.15 0.87 0.365 0.8 0.365 0.8 0.22 0.495 0.22 0.495 0.5 0.045 0.5  ;
  END
END OAI22_X1

MACRO OAI22_X2
  CLASS core ;
  FOREIGN OAI22_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.065 1.315 0.065 1.065 0.135 1.065 0.135 1.315 0.82 1.315 0.82 1.065 0.89 1.065 0.89 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.56 0.375 0.56 0.375 0.7 0.25 0.7  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.56 0.565 0.56 0.565 0.7 0.44 0.7  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.32 0.085 0.32 0.235 0.25 0.235 0.25 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.185 0.56 0.185 0.7 0.06 0.7  ;
    END
  END B2
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.765 0.42 0.89 0.42 0.89 0.56 0.765 0.56  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.45 0.765 0.63 0.765 0.63 0.285 0.7 0.285 0.7 0.835 0.52 0.835 0.52 1.165 0.45 1.165  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.035 0.3 0.44 0.3 0.44 0.15 0.89 0.15 0.89 0.285 0.82 0.285 0.82 0.22 0.51 0.22 0.51 0.37 0.035 0.37  ;
  END
END OAI22_X2

MACRO OAI22_X4
  CLASS core ;
  FOREIGN OAI22_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.71 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 1.065 0.115 1.065 0.115 1.315 0.77 1.315 0.77 1.1 0.905 1.1 0.905 1.315 1.56 1.315 1.56 1.065 1.63 1.065 1.63 1.315 1.71 1.315 1.71 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.7 0.41 0.7 0.41 0.84 0.25 0.84  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.2 0.76 1.335 0.76 1.335 0.98 1.2 0.98  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.71 -0.085 1.71 0.085 0.72 0.085 0.72 0.205 0.585 0.205 0.585 0.085 0.34 0.085 0.34 0.205 0.205 0.205 0.205 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.12 0.56 0.755 0.56 0.755 0.7 0.63 0.7 0.63 0.63 0.12 0.63  ;
    END
  END B2
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.955 0.56 1.56 0.56 1.56 0.63 1.08 0.63 1.08 0.7 0.955 0.7  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.43 0.91 0.82 0.91 0.82 0.425 0.96 0.425 0.96 0.325 1.475 0.325 1.475 0.395 1.03 0.395 1.03 0.495 0.89 0.495 0.89 0.91 1.07 0.91 1.07 1.045 1.285 1.045 1.285 1.115 1 1.115 1 0.98 0.5 0.98 0.5 1.185 0.43 1.185  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.05 0.225 0.12 0.225 0.12 0.29 0.8 0.29 0.8 0.15 1.63 0.15 1.63 0.425 1.56 0.425 1.56 0.22 0.87 0.22 0.87 0.36 0.05 0.36  ;
  END
END OAI22_X4

MACRO OAI33_X1
  CLASS core ;
  FOREIGN OAI33_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.33 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.055 1.315 0.055 1.065 0.125 1.065 0.125 1.315 1.19 1.315 1.19 1.065 1.26 1.065 1.26 1.315 1.33 1.315 1.33 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.98 0.495 0.98 0.495 0.675 0.565 0.675 0.565 1.12 0.44 1.12  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.765 0.7 0.89 0.7 0.89 0.84 0.765 0.84  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.955 0.84 1.08 0.84 1.08 0.98 0.955 0.98  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 0.565 0.81 0.565 0.81 0.285 0.88 0.285 0.88 0.565 1.19 0.565 1.19 0.285 1.26 0.285 1.26 0.635 0.7 0.635 0.7 1.155 0.63 1.155  ;
    END
  END ZN
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.145 0.84 1.27 0.84 1.27 0.98 1.145 0.98  ;
    END
  END A3
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.185 0.56 0.185 0.7 0.06 0.7  ;
    END
  END B3
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.33 -0.085 1.33 0.085 0.5 0.085 0.5 0.365 0.43 0.365 0.43 0.085 0.125 0.085 0.125 0.365 0.055 0.365 0.055 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.78 0.42 0.78 0.42 0.915 0.32 0.915 0.32 0.98 0.25 0.98  ;
    END
  END B2
  OBS
      LAYER metal1 ;
        POLYGON 0.25 0.285 0.32 0.285 0.32 0.43 0.63 0.43 0.63 0.15 1.07 0.15 1.07 0.365 1 0.365 1 0.22 0.7 0.22 0.7 0.5 0.25 0.5  ;
  END
END OAI33_X1

MACRO OR2_X1
  CLASS core ;
  FOREIGN OR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.42 1.315 0.42 1.145 0.49 1.145 0.49 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.17 0.925 0.245 0.925 0.245 1.155 0.355 1.155 0.355 1.225 0.175 1.225 0.175 1.06 0.17 1.06  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.485 0.085 0.485 0.27 0.415 0.27 0.415 0.085 0.11 0.085 0.11 0.27 0.04 0.27 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.315 0.56 0.51 0.56 0.51 0.7 0.315 0.7  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 0.15 0.7 0.15 0.7 1.22 0.63 1.22  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.035 0.335 0.225 0.335 0.225 0.15 0.295 0.15 0.295 0.335 0.565 0.335 0.565 0.405 0.105 0.405 0.105 1.085 0.11 1.085 0.11 1.22 0.035 1.22  ;
  END
END OR2_X1

MACRO OR2_X2
  CLASS core ;
  FOREIGN OR2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.415 1.315 0.415 1.17 0.485 1.17 0.485 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.17 0.42 0.17 0.56 0.06 0.56  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.51 0.085 0.51 0.195 0.44 0.195 0.44 0.085 0.11 0.085 0.11 0.285 0.04 0.285 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.37 0.56 0.51 0.56 0.51 0.7 0.37 0.7  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 0.165 0.7 0.165 0.7 1.25 0.63 1.25  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.625 0.235 0.625 0.235 0.165 0.305 0.165 0.305 0.425 0.565 0.425 0.565 0.495 0.305 0.495 0.305 0.695 0.115 0.695 0.115 1.185 0.045 1.185  ;
  END
END OR2_X2

MACRO OR2_X4
  CLASS core ;
  FOREIGN OR2_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.425 1.315 0.425 1.205 0.495 1.205 0.495 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.15 0.42 0.15 0.56 0.06 0.56  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.495 0.085 0.495 0.27 0.425 0.27 0.425 0.085 0.12 0.085 0.12 0.27 0.05 0.27 0.05 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.35 0.455 0.545 0.455 0.545 0.525 0.42 0.525 0.42 0.655 0.35 0.655  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 0.28 0.7 0.28 0.7 1.015 0.63 1.015  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.285 0.735 0.495 0.735 0.495 0.615 0.565 0.615 0.565 0.805 0.125 0.805 0.125 1.22 0.055 1.22 0.055 0.735 0.215 0.735 0.215 0.15 0.305 0.15 0.305 0.285 0.285 0.285  ;
  END
END OR2_X4

MACRO OR3_X1
  CLASS core ;
  FOREIGN OR3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.64 1.315 0.64 1.035 0.71 1.035 0.71 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.505 0.875 0.735 0.875 0.735 0.945 0.505 0.945  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.185 0.56 0.32 0.56 0.32 0.7 0.185 0.7  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.71 0.085 0.71 0.27 0.64 0.27 0.64 0.085 0.33 0.085 0.33 0.27 0.26 0.27 0.26 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.385 0.56 0.51 0.56 0.51 0.7 0.385 0.7  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.82 0.15 0.9 0.15 0.9 1.11 0.82 1.11  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.05 0.15 0.145 0.15 0.145 0.335 0.45 0.335 0.45 0.15 0.52 0.15 0.52 0.335 0.755 0.335 0.755 0.47 0.685 0.47 0.685 0.405 0.12 0.405 0.12 0.975 0.145 0.975 0.145 1.25 0.05 1.25  ;
  END
END OR3_X1

MACRO OR3_X2
  CLASS core ;
  FOREIGN OR3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.63 1.315 0.63 1.205 0.7 1.205 0.7 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.53 0.895 0.7 0.895 0.7 1.12 0.63 1.12 0.63 1.03 0.53 1.03  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.175 0.56 0.32 0.56 0.32 0.7 0.175 0.7  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.7 0.085 0.7 0.27 0.63 0.27 0.63 0.085 0.32 0.085 0.32 0.27 0.25 0.27 0.25 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.385 0.56 0.51 0.56 0.51 0.7 0.385 0.7  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.82 0.24 0.89 0.24 0.89 1.145 0.82 1.145  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.04 0.15 0.135 0.15 0.135 0.365 0.445 0.365 0.445 0.15 0.525 0.15 0.525 0.365 0.755 0.365 0.755 0.5 0.685 0.5 0.685 0.435 0.11 0.435 0.11 1.02 0.135 1.02 0.135 1.155 0.04 1.155  ;
  END
END OR3_X2

MACRO OR3_X4
  CLASS core ;
  FOREIGN OR3_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.625 1.315 0.625 0.925 0.695 0.925 0.695 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.525 0.615 0.595 0.615 0.595 0.7 0.7 0.7 0.7 0.84 0.525 0.84  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.98 0.195 0.98 0.195 0.715 0.19 0.715 0.19 0.58 0.265 0.58 0.265 1.12 0.06 1.12  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.695 0.085 0.695 0.27 0.625 0.27 0.625 0.085 0.315 0.085 0.315 0.27 0.245 0.27 0.245 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.36 0.615 0.43 0.615 0.43 0.98 0.51 0.98 0.51 1.12 0.36 1.12  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.82 0.205 0.89 0.205 0.89 1.015 0.82 1.015  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.055 0.15 0.13 0.15 0.13 0.335 0.435 0.335 0.435 0.15 0.505 0.15 0.505 0.335 0.755 0.335 0.755 0.605 0.685 0.605 0.685 0.405 0.125 0.405 0.125 0.74 0.13 0.74 0.13 0.875 0.055 0.875  ;
  END
END OR3_X4

MACRO OR4_X1
  CLASS core ;
  FOREIGN OR4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.82 1.315 0.82 1.015 0.89 1.015 0.89 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.575 0.56 0.7 0.56 0.7 0.7 0.575 0.7  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.175 0.56 0.32 0.56 0.32 0.7 0.175 0.7  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.89 0.085 0.89 0.27 0.82 0.27 0.82 0.085 0.51 0.085 0.51 0.27 0.44 0.27 0.44 0.085 0.135 0.085 0.135 0.27 0.065 0.27 0.065 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.385 0.7 0.51 0.7 0.51 0.84 0.385 0.84  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.765 0.56 0.89 0.56 0.89 0.7 0.765 0.7  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.01 0.98 1.035 0.98 1.035 0.285 1.015 0.285 1.015 0.15 1.105 0.15 1.105 1.12 1.01 1.12  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.04 0.335 0.25 0.335 0.25 0.15 0.32 0.15 0.32 0.335 0.63 0.335 0.63 0.15 0.7 0.15 0.7 0.335 0.97 0.335 0.97 0.405 0.11 0.405 0.11 0.955 0.135 0.955 0.135 1.23 0.04 1.23  ;
  END
END OR4_X1

MACRO OR4_X2
  CLASS core ;
  FOREIGN OR4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.815 1.315 0.815 1.01 0.885 1.01 0.885 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.575 0.56 0.7 0.56 0.7 0.7 0.575 0.7  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.17 0.56 0.32 0.56 0.32 0.7 0.17 0.7  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.885 0.085 0.885 0.27 0.815 0.27 0.815 0.085 0.505 0.085 0.505 0.27 0.435 0.27 0.435 0.085 0.13 0.085 0.13 0.27 0.06 0.27 0.06 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.385 0.56 0.51 0.56 0.51 0.7 0.385 0.7  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.765 0.56 0.89 0.56 0.89 0.7 0.765 0.7  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.01 0.56 1.03 0.56 1.03 0.22 1.1 0.22 1.1 1.09 1.01 1.09  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.035 0.375 0.245 0.375 0.245 0.15 0.315 0.15 0.315 0.375 0.625 0.375 0.625 0.15 0.695 0.15 0.695 0.375 0.965 0.375 0.965 0.445 0.105 0.445 0.105 0.955 0.13 0.955 0.13 1.23 0.035 1.23  ;
  END
END OR4_X2

MACRO OR4_X4
  CLASS core ;
  FOREIGN OR4_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.815 1.315 0.815 1.065 0.885 1.065 0.885 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.405 0.455 0.55 0.455 0.55 0.59 0.405 0.59  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.18 0.42 0.18 0.56 0.06 0.56  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.885 0.085 0.885 0.27 0.815 0.27 0.815 0.085 0.54 0.085 0.54 0.235 0.405 0.235 0.405 0.085 0.13 0.085 0.13 0.27 0.06 0.27 0.06 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.38 0.7 0.51 0.7 0.51 0.84 0.38 0.84  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.715 0.695 0.89 0.695 0.89 0.84 0.715 0.84  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.01 0.165 1.08 0.165 1.08 1.155 1.01 1.155  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.065 0.925 0.245 0.925 0.245 0.15 0.315 0.15 0.315 0.315 0.625 0.315 0.625 0.15 0.695 0.15 0.695 0.43 0.945 0.43 0.945 0.565 0.625 0.565 0.625 0.385 0.315 0.385 0.315 0.995 0.135 0.995 0.135 1.23 0.065 1.23  ;
  END
END OR4_X4

MACRO SDFFRS_X1
  CLASS core ;
  FOREIGN SDFFRS_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 6.27 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 5.74 0.405 5.83 0.405 5.83 0.915 5.74 0.915  ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.885 0.68 4.79 0.68 4.79 0.815 4.585 0.815 4.585 0.75 2.885 0.75  ;
    END
  END SN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.18 0.815 0.32 0.815 0.32 0.98 0.18 0.98  ;
    END
  END SE
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 5.19 0.42 5.375 0.42 5.375 0.56 5.19 0.56  ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.265 1.315 0.265 1.2 0.4 1.2 0.4 1.315 1.02 1.315 1.02 1.2 1.155 1.2 1.155 1.315 1.41 1.315 1.41 0.95 1.545 0.95 1.545 1.315 2.215 1.315 2.215 1.115 2.35 1.115 2.35 1.315 2.99 1.315 2.99 1.115 3.125 1.115 3.125 1.315 3.55 1.315 3.55 1.115 3.685 1.115 3.685 1.315 4.105 1.315 4.105 1.19 4.24 1.19 4.24 1.315 4.95 1.315 4.95 1.19 5.085 1.19 5.085 1.315 5.365 1.315 5.365 1.115 5.5 1.115 5.5 1.315 5.74 1.315 5.74 1.16 5.925 1.16 5.925 0.84 5.995 0.84 5.995 1.315 6.27 1.315 6.27 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 6.115 0.28 6.21 0.28 6.21 0.915 6.115 0.915  ;
    END
  END Q
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.42 0.46 0.42 0.46 0.56 0.25 0.56  ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 5.895 0.42 5.98 0.42 5.98 0.085 5.33 0.085 5.33 0.21 5.195 0.21 5.195 0.085 4.72 0.085 4.72 0.285 4.585 0.285 4.585 0.085 3.67 0.085 3.67 0.285 3.535 0.285 3.535 0.085 2.955 0.085 2.955 0.34 2.82 0.34 2.82 0.085 1.925 0.085 1.925 0.34 1.79 0.34 1.79 0.085 1.55 0.085 1.55 0.21 1.415 0.21 1.415 0.085 1.135 0.085 1.135 0.285 1 0.285 1 0.085 0.38 0.085 0.38 0.285 0.245 0.285 0.245 0.085 0 0.085 0 -0.085 6.27 -0.085 6.27 0.085 6.05 0.085 6.05 0.49 5.895 0.49  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.385 0.78 0.93 0.78 0.93 0.485 1 0.485 1 0.85 0.52 0.85 0.52 0.98 0.385 0.98  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.37 0.34 1.39 0.34 1.39 0.28 1.46 0.28 1.46 0.475 1.37 0.475  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.29 0.14 0.29 0.14 0.645 0.865 0.645 0.865 0.715 0.115 0.715 0.115 1.18 0.2 1.18 0.2 1.25 0.045 1.25  ;
        POLYGON 1.295 0.565 1.63 0.565 1.63 0.635 1.36 0.635 1.36 0.73 1.225 0.73 1.225 0.155 1.325 0.155 1.325 0.29 1.295 0.29  ;
        POLYGON 3.765 1.055 4.185 1.055 4.185 0.815 4.255 0.815 4.255 1.055 5.02 1.055 5.02 0.78 5.39 0.78 5.39 0.85 5.09 0.85 5.09 1.125 4.71 1.125 4.71 1.195 4.575 1.195 4.575 1.125 3.835 1.125 3.835 1.23 3.765 1.23  ;
        POLYGON 5.155 0.915 5.47 0.915 5.47 0.355 5.095 0.355 5.095 0.425 4.35 0.425 4.35 0.35 5.025 0.35 5.025 0.285 5.54 0.285 5.54 0.985 5.155 0.985  ;
        POLYGON 5.59 1.065 5.605 1.065 5.605 0.165 5.915 0.165 5.915 0.24 5.675 0.24 5.675 1.2 5.59 1.2  ;
        POLYGON 0.645 0.915 1.065 0.915 1.065 0.42 0.625 0.42 0.625 0.325 0.76 0.325 0.76 0.35 1.135 0.35 1.135 0.8 1.8 0.8 1.8 0.705 1.87 0.705 1.87 0.87 1.135 0.87 1.135 0.985 0.645 0.985  ;
        POLYGON 2.21 0.15 2.345 0.15 2.345 0.355 2.21 0.355  ;
        POLYGON 2.095 0.555 2.165 0.555 2.165 0.805 2.745 0.805 2.745 1 2.61 1 2.61 0.875 2.095 0.875  ;
        POLYGON 2.55 0.41 3.02 0.41 3.02 0.235 3.155 0.235 3.155 0.41 3.385 0.41 3.385 0.48 2.55 0.48  ;
        POLYGON 3.225 0.95 3.36 0.95 3.36 1.055 3.485 1.055 3.485 1.125 3.225 1.125  ;
        POLYGON 1.805 1.095 2.075 1.095 2.075 0.965 2.49 0.965 2.49 1.095 2.855 1.095 2.855 0.815 4.12 0.815 4.12 0.99 3.985 0.99 3.985 0.885 2.925 0.885 2.925 1.165 2.42 1.165 2.42 1.035 2.145 1.035 2.145 1.165 1.805 1.165  ;
        POLYGON 3.955 0.185 4.045 0.185 4.045 0.41 4.285 0.41 4.285 0.48 3.975 0.48 3.975 0.32 3.955 0.32  ;
        POLYGON 4.655 0.92 4.855 0.92 4.855 0.615 2.415 0.615 2.415 0.49 2.01 0.49 2.01 1.03 1.61 1.03 1.61 0.95 1.94 0.95 1.94 0.49 1.635 0.49 1.635 0.215 1.705 0.215 1.705 0.42 2.485 0.42 2.485 0.545 3.84 0.545 3.84 0.37 3.91 0.37 3.91 0.545 4.925 0.545 4.925 0.99 4.655 0.99  ;
  END
END SDFFRS_X1

MACRO SDFFRS_X2
  CLASS core ;
  FOREIGN SDFFRS_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 6.27 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 5.74 0.405 5.83 0.405 5.83 0.56 5.81 0.56 5.81 0.915 5.74 0.915  ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.885 0.68 4.79 0.68 4.79 0.815 4.585 0.815 4.585 0.75 2.885 0.75  ;
    END
  END SN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.18 0.815 0.32 0.815 0.32 0.98 0.18 0.98  ;
    END
  END SE
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 5.19 0.42 5.375 0.42 5.375 0.56 5.19 0.56  ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.265 1.315 0.265 1.2 0.4 1.2 0.4 1.315 1.02 1.315 1.02 1.2 1.155 1.2 1.155 1.315 1.41 1.315 1.41 0.95 1.545 0.95 1.545 1.315 2.215 1.315 2.215 1.23 2.35 1.23 2.35 1.315 2.99 1.315 2.99 1.115 3.125 1.115 3.125 1.315 3.55 1.315 3.55 1.115 3.685 1.115 3.685 1.315 4.105 1.315 4.105 1.19 4.24 1.19 4.24 1.315 4.95 1.315 4.95 1.19 5.085 1.19 5.085 1.315 5.365 1.315 5.365 1.115 5.5 1.115 5.5 1.315 5.74 1.315 5.74 1.16 5.89 1.16 5.89 0.875 6.025 0.875 6.025 1.315 6.27 1.315 6.27 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 6.115 0.28 6.21 0.28 6.21 0.915 6.115 0.915  ;
    END
  END Q
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.42 0.46 0.42 0.46 0.56 0.25 0.56  ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 5.895 0.42 5.98 0.42 5.98 0.085 5.23 0.085 5.23 0.21 5.095 0.21 5.095 0.085 4.72 0.085 4.72 0.285 4.585 0.285 4.585 0.085 3.67 0.085 3.67 0.285 3.535 0.285 3.535 0.085 2.955 0.085 2.955 0.34 2.82 0.34 2.82 0.085 1.925 0.085 1.925 0.34 1.79 0.34 1.79 0.085 1.55 0.085 1.55 0.21 1.415 0.21 1.415 0.085 1.135 0.085 1.135 0.285 1 0.285 1 0.085 0.38 0.085 0.38 0.285 0.245 0.285 0.245 0.085 0 0.085 0 -0.085 6.27 -0.085 6.27 0.085 6.05 0.085 6.05 0.49 5.895 0.49  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.385 0.78 0.93 0.78 0.93 0.485 1 0.485 1 0.85 0.52 0.85 0.52 0.98 0.385 0.98  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.37 0.34 1.39 0.34 1.39 0.28 1.46 0.28 1.46 0.475 1.37 0.475  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.29 0.14 0.29 0.14 0.645 0.865 0.645 0.865 0.715 0.115 0.715 0.115 1.18 0.2 1.18 0.2 1.25 0.045 1.25  ;
        POLYGON 1.295 0.66 1.655 0.66 1.655 0.73 1.225 0.73 1.225 0.155 1.325 0.155 1.325 0.29 1.295 0.29  ;
        POLYGON 3.765 1.055 4.185 1.055 4.185 0.815 4.255 0.815 4.255 1.055 5.02 1.055 5.02 0.78 5.39 0.78 5.39 0.85 5.09 0.85 5.09 1.125 4.71 1.125 4.71 1.195 4.575 1.195 4.575 1.125 3.835 1.125 3.835 1.23 3.765 1.23  ;
        POLYGON 5.155 0.915 5.47 0.915 5.47 0.355 5.095 0.355 5.095 0.425 4.35 0.425 4.35 0.35 5.025 0.35 5.025 0.285 5.54 0.285 5.54 0.985 5.155 0.985  ;
        POLYGON 5.59 1.065 5.605 1.065 5.605 0.22 5.52 0.22 5.52 0.15 5.795 0.15 5.795 0.22 5.675 0.22 5.675 1.2 5.59 1.2  ;
        POLYGON 0.645 0.915 1.065 0.915 1.065 0.42 0.625 0.42 0.625 0.325 0.76 0.325 0.76 0.35 1.135 0.35 1.135 0.81 1.8 0.81 1.8 0.725 1.87 0.725 1.87 0.88 1.135 0.88 1.135 0.985 0.645 0.985  ;
        POLYGON 2.21 0.15 2.345 0.15 2.345 0.355 2.21 0.355  ;
        POLYGON 2.095 0.555 2.165 0.555 2.165 0.96 2.665 0.96 2.665 1.03 2.095 1.03  ;
        POLYGON 2.55 0.41 3.02 0.41 3.02 0.235 3.155 0.235 3.155 0.41 3.385 0.41 3.385 0.48 2.55 0.48  ;
        POLYGON 3.225 0.95 3.36 0.95 3.36 1.055 3.485 1.055 3.485 1.125 3.225 1.125  ;
        POLYGON 1.805 1.095 2.855 1.095 2.855 0.815 4.12 0.815 4.12 0.99 3.985 0.99 3.985 0.885 2.925 0.885 2.925 1.17 2.61 1.17 2.61 1.165 1.805 1.165  ;
        POLYGON 3.955 0.185 4.045 0.185 4.045 0.41 4.285 0.41 4.285 0.48 3.975 0.48 3.975 0.32 3.955 0.32  ;
        POLYGON 4.655 0.92 4.855 0.92 4.855 0.615 2.415 0.615 2.415 0.49 2.01 0.49 2.01 1.03 1.61 1.03 1.61 0.95 1.94 0.95 1.94 0.49 1.635 0.49 1.635 0.215 1.705 0.215 1.705 0.42 2.485 0.42 2.485 0.545 3.84 0.545 3.84 0.37 3.91 0.37 3.91 0.545 4.925 0.545 4.925 0.99 4.655 0.99  ;
  END
END SDFFRS_X2

MACRO SDFFR_X1
  CLASS core ;
  FOREIGN SDFFR_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 4.94 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.05 0.15 0.13 0.15 0.13 0.95 0.05 0.95  ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 4.24 0.56 4.34 0.56 4.34 0.7 4.24 0.7  ;
    END
  END SE
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.355 0.81 2.645 0.81 2.645 0.88 1.495 0.88 1.495 0.945 1.355 0.945  ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.23 1.315 0.23 0.875 0.3 0.875 0.3 1.315 0.735 1.315 0.735 1.115 0.805 1.115 0.805 1.315 1.485 1.315 1.485 1.28 1.62 1.28 1.62 1.315 2.265 1.315 2.265 0.995 2.335 0.995 2.335 1.315 2.645 1.315 2.645 1.13 2.715 1.13 2.715 1.315 3.42 1.315 3.42 0.995 3.49 0.995 3.49 1.315 3.81 1.315 3.81 1.065 3.88 1.065 3.88 1.315 4.57 1.315 4.57 1.065 4.64 1.065 4.64 1.315 4.94 1.315 4.94 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.42 0.15 0.51 0.15 0.51 0.42 0.49 0.42 0.49 0.95 0.42 0.95  ;
    END
  END Q
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 4.43 0.52 4.53 0.52 4.53 0.7 4.43 0.7  ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 4.94 -0.085 4.94 0.085 4.635 0.085 4.635 0.32 4.565 0.32 4.565 0.085 3.88 0.085 3.88 0.32 3.81 0.32 3.81 0.085 3.465 0.085 3.465 0.235 3.395 0.235 3.395 0.085 2.725 0.085 2.725 0.2 2.59 0.2 2.59 0.085 1.78 0.085 1.78 0.235 1.71 0.235 1.71 0.085 0.835 0.085 0.835 0.235 0.765 0.235 0.765 0.085 0.305 0.085 0.305 0.27 0.235 0.27 0.235 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.92 0.53 3.995 0.53 3.995 0.795 4.53 0.795 4.53 1.01 4.5 1.01 4.5 1.12 4.43 1.12 4.43 0.865 3.92 0.865  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.445 0.595 3.61 0.595 3.61 0.665 3.445 0.665  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.555 0.6 0.575 0.6 0.575 0.155 0.645 0.155 0.645 0.67 0.625 0.67 0.625 1.235 0.555 1.235  ;
        POLYGON 1.055 1.145 2.03 1.145 2.03 1.215 0.985 1.215 0.985 1.05 0.69 1.05 0.69 0.915 0.71 0.915 0.71 0.42 0.78 0.42 0.78 0.98 0.985 0.98 0.985 0.15 1.435 0.15 1.435 0.22 1.055 0.22  ;
        POLYGON 2.43 0.995 2.745 0.995 2.745 0.81 2.815 0.81 2.815 1.065 2.565 1.065 2.565 1.08 2.43 1.08  ;
        POLYGON 2.215 0.15 2.35 0.15 2.35 0.27 2.835 0.27 2.835 0.34 2.215 0.34  ;
        POLYGON 1.12 0.3 1.9 0.3 1.9 0.205 1.97 0.205 1.97 0.405 2.9 0.405 2.9 0.34 2.97 0.34 2.97 0.475 1.9 0.475 1.9 0.435 1.19 0.435 1.19 1.01 2.185 1.01 2.185 1.08 1.12 1.08  ;
        POLYGON 1.6 0.54 3.035 0.54 3.035 0.305 3.025 0.305 3.025 0.17 3.105 0.17 3.105 0.54 3.115 0.54 3.115 1.115 3.045 1.115 3.045 0.61 1.6 0.61  ;
        POLYGON 3.25 0.86 3.68 0.86 3.68 1.025 3.61 1.025 3.61 0.93 3.25 0.93 3.25 1.25 2.91 1.25 2.91 0.745 1.255 0.745 1.255 0.5 1.325 0.5 1.325 0.675 2.98 0.675 2.98 1.18 3.18 1.18 3.18 0.465 3.17 0.465 3.17 0.3 3.585 0.3 3.585 0.205 3.655 0.205 3.655 0.37 3.25 0.37  ;
        POLYGON 3.315 0.435 3.785 0.435 3.785 0.395 3.97 0.395 3.97 0.25 4.29 0.25 4.29 0.32 4.04 0.32 4.04 0.465 3.855 0.465 3.855 0.93 4.255 0.93 4.255 1.145 4.185 1.145 4.185 1 3.785 1 3.785 0.505 3.385 0.505 3.385 0.57 3.315 0.57  ;
        POLYGON 4.105 0.385 4.755 0.385 4.755 0.29 4.825 0.29 4.825 1.145 4.755 1.145 4.755 0.455 4.175 0.455 4.175 0.55 4.105 0.55  ;
  END
END SDFFR_X1

MACRO SDFFR_X2
  CLASS core ;
  FOREIGN SDFFR_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 4.94 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.05 0.165 0.13 0.165 0.13 0.915 0.05 0.915  ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 4.24 0.56 4.335 0.56 4.335 0.7 4.24 0.7  ;
    END
  END SE
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.355 0.81 2.625 0.81 2.625 0.88 1.495 0.88 1.495 0.945 1.355 0.945  ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.23 1.315 0.23 0.975 0.3 0.975 0.3 1.315 0.74 1.315 0.74 1.13 0.81 1.13 0.81 1.315 1.485 1.315 1.485 1.28 1.62 1.28 1.62 1.315 2.265 1.315 2.265 0.995 2.335 0.995 2.335 1.315 2.615 1.315 2.615 1.165 2.75 1.165 2.75 1.315 3.42 1.315 3.42 0.995 3.49 0.995 3.49 1.315 3.805 1.315 3.805 1.065 3.875 1.065 3.875 1.315 4.565 1.315 4.565 1.205 4.635 1.205 4.635 1.315 4.94 1.315 4.94 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.42 0.165 0.51 0.165 0.51 0.42 0.49 0.42 0.49 0.915 0.42 0.915  ;
    END
  END Q
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 4.43 0.52 4.525 0.52 4.525 0.7 4.43 0.7  ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 4.94 -0.085 4.94 0.085 4.63 0.085 4.63 0.32 4.56 0.32 4.56 0.085 3.88 0.085 3.88 0.32 3.81 0.32 3.81 0.085 3.445 0.085 3.445 0.195 3.375 0.195 3.375 0.085 2.705 0.085 2.705 0.16 2.57 0.16 2.57 0.085 1.78 0.085 1.78 0.285 1.71 0.285 1.71 0.085 0.84 0.085 0.84 0.285 0.77 0.285 0.77 0.085 0.305 0.085 0.305 0.195 0.235 0.195 0.235 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.915 0.53 3.985 0.53 3.985 0.795 4.525 0.795 4.525 1.12 4.43 1.12 4.43 0.865 3.915 0.865  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.435 0.56 3.555 0.56 3.555 0.7 3.435 0.7  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.555 0.53 0.575 0.53 0.575 0.255 0.645 0.255 0.645 0.6 0.625 0.6 0.625 1.25 0.555 1.25  ;
        POLYGON 1.03 1.145 2.03 1.145 2.03 1.215 0.96 1.215 0.96 0.45 0.78 0.45 0.78 0.815 0.7 0.815 0.7 0.68 0.71 0.68 0.71 0.38 0.96 0.38 0.96 0.2 1.435 0.2 1.435 0.27 1.03 0.27  ;
        POLYGON 2.43 1.01 2.735 1.01 2.735 0.855 2.805 0.855 2.805 1.08 2.43 1.08  ;
        POLYGON 2.175 0.15 2.31 0.15 2.31 0.25 2.815 0.25 2.815 0.32 2.175 0.32  ;
        POLYGON 1.095 0.385 1.9 0.385 1.9 0.165 1.97 0.165 1.97 0.385 2.88 0.385 2.88 0.32 2.95 0.32 2.95 0.455 1.165 0.455 1.165 1.01 2.185 1.01 2.185 1.08 1.095 1.08  ;
        POLYGON 1.6 0.54 3.015 0.54 3.015 0.285 3.005 0.285 3.005 0.15 3.085 0.15 3.085 0.98 3.11 0.98 3.11 1.115 3.015 1.115 3.015 0.61 1.6 0.61  ;
        POLYGON 3.22 0.83 3.715 0.83 3.715 0.9 3.245 0.9 3.245 1.25 2.88 1.25 2.88 0.745 1.23 0.745 1.23 0.52 1.3 0.52 1.3 0.675 2.95 0.675 2.95 1.18 3.175 1.18 3.175 0.9 3.15 0.9 3.15 0.26 3.565 0.26 3.565 0.165 3.635 0.165 3.635 0.33 3.22 0.33  ;
        POLYGON 3.285 0.395 3.97 0.395 3.97 0.25 4.285 0.25 4.285 0.32 4.04 0.32 4.04 0.465 3.85 0.465 3.85 0.93 4.25 0.93 4.25 1.145 4.18 1.145 4.18 1 3.78 1 3.78 0.465 3.285 0.465  ;
        POLYGON 4.105 0.385 4.75 0.385 4.75 0.29 4.82 0.29 4.82 1.145 4.75 1.145 4.75 0.455 4.175 0.455 4.175 0.55 4.105 0.55  ;
  END
END SDFFR_X2

MACRO SDFFS_X1
  CLASS core ;
  FOREIGN SDFFS_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 5.13 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 4.585 0.15 4.655 0.15 4.655 0.28 4.69 0.28 4.69 0.42 4.655 0.42 4.655 1.155 4.585 1.155  ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.67 0.275 3.93 0.275 3.93 0.53 4.19 0.53 4.19 0.6 3.86 0.6 3.86 0.345 2.74 0.345 2.74 0.46 2.67 0.46  ;
    END
  END SN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.22 0.42 0.32 0.42 0.32 0.7 0.22 0.7  ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.265 1.315 0.265 1.24 0.4 1.24 0.4 1.315 1.025 1.315 1.025 1.24 1.16 1.24 1.16 1.315 1.76 1.315 1.76 1.095 1.41 1.095 1.41 1.025 1.83 1.025 1.83 1.315 2.485 1.315 2.485 1.1 2.62 1.1 2.62 1.315 3.04 1.315 3.04 1.115 3.175 1.115 3.175 1.315 3.95 1.315 3.95 1.115 4.085 1.115 4.085 1.315 4.34 1.315 4.34 1.115 4.475 1.115 4.475 1.315 4.765 1.315 4.765 1.08 4.835 1.08 4.835 1.315 5.13 1.315 5.13 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 4.96 0.15 5.07 0.15 5.07 1.155 4.96 1.155  ;
    END
  END Q
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.385 0.415 0.51 0.415 0.51 0.56 0.385 0.56  ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 5.13 -0.085 5.13 0.085 4.875 0.085 4.875 0.235 4.74 0.235 4.74 0.085 4.13 0.085 4.13 0.42 3.995 0.42 3.995 0.085 2.895 0.085 2.895 0.21 2.76 0.21 2.76 0.085 1.9 0.085 1.9 0.32 1.83 0.32 1.83 0.085 1.55 0.085 1.55 0.21 1.415 0.21 1.415 0.085 1.135 0.085 1.135 0.285 1 0.285 1 0.085 0.34 0.085 0.34 0.32 0.27 0.32 0.27 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.375 0.92 0.93 0.92 0.93 0.485 1 0.485 1 0.99 0.51 0.99 0.51 1.12 0.375 1.12  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.39 0.56 1.475 0.56 1.475 0.7 1.39 0.7  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.085 0.29 0.155 0.29 0.155 0.785 0.865 0.785 0.865 0.855 0.18 0.855 0.18 1.145 0.085 1.145  ;
        POLYGON 1.295 0.415 1.63 0.415 1.63 0.485 1.295 0.485 1.295 0.83 1.36 0.83 1.36 0.9 1.225 0.9 1.225 0.25 1.36 0.25 1.36 0.32 1.295 0.32  ;
        POLYGON 0.65 1.055 1.065 1.055 1.065 0.42 0.625 0.42 0.625 0.325 0.76 0.325 0.76 0.35 1.135 0.35 1.135 1.055 1.295 1.055 1.295 1.18 1.695 1.18 1.695 1.25 1.225 1.25 1.225 1.125 0.65 1.125  ;
        POLYGON 1.65 0.795 1.695 0.795 1.695 0.35 1.635 0.35 1.635 0.215 1.765 0.215 1.765 0.675 2.11 0.675 2.11 0.745 1.765 0.745 1.765 0.93 1.65 0.93  ;
        POLYGON 2.065 0.45 2.245 0.45 2.245 0.905 2.175 0.905 2.175 0.52 2.065 0.52  ;
        POLYGON 2.445 0.525 2.955 0.525 2.955 0.44 3.09 0.44 3.09 0.645 3.175 0.645 3.175 0.715 3.02 0.715 3.02 0.595 2.445 0.595  ;
        POLYGON 2.14 0.97 2.31 0.97 2.31 0.305 2.175 0.305 2.175 0.235 2.38 0.235 2.38 0.81 3.255 0.81 3.255 0.73 3.325 0.73 3.325 0.88 2.38 0.88 2.38 1.04 2.21 1.04 2.21 1.185 2.14 1.185  ;
        POLYGON 3.375 0.41 3.445 0.41 3.445 0.545 3.66 0.545 3.66 0.895 3.59 0.895 3.59 0.615 3.375 0.615  ;
        POLYGON 3.515 0.96 3.725 0.96 3.725 0.48 3.51 0.48 3.51 0.41 3.795 0.41 3.795 0.78 4.37 0.78 4.37 0.85 3.795 0.85 3.795 1.03 3.515 1.03  ;
        POLYGON 3.86 0.915 4.45 0.915 4.45 0.51 4.405 0.51 4.405 0.235 4.52 0.235 4.52 0.985 3.86 0.985  ;
  END
END SDFFS_X1

MACRO SDFFS_X2
  CLASS core ;
  FOREIGN SDFFS_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 5.13 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 4.585 0.15 4.655 0.15 4.655 0.42 4.69 0.42 4.69 0.56 4.655 0.56 4.655 1.02 4.585 1.02  ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.67 0.275 3.93 0.275 3.93 0.53 4.19 0.53 4.19 0.6 3.86 0.6 3.86 0.345 2.74 0.345 2.74 0.46 2.67 0.46  ;
    END
  END SN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.22 0.42 0.32 0.42 0.32 0.7 0.22 0.7  ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.265 1.315 0.265 1.24 0.4 1.24 0.4 1.315 1.025 1.315 1.025 1.24 1.16 1.24 1.16 1.315 1.76 1.315 1.76 1.095 1.41 1.095 1.41 1.025 1.83 1.025 1.83 1.315 2.485 1.315 2.485 1.1 2.62 1.1 2.62 1.315 3.04 1.315 3.04 1.115 3.175 1.115 3.175 1.315 3.95 1.315 3.95 1.115 4.085 1.115 4.085 1.315 4.34 1.315 4.34 1.115 4.475 1.115 4.475 1.315 4.765 1.315 4.765 1.08 4.835 1.08 4.835 1.315 5.13 1.315 5.13 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 4.96 0.885 5 0.885 5 0.345 4.96 0.345 4.96 0.15 5.07 0.15 5.07 1.02 4.96 1.02  ;
    END
  END Q
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.385 0.415 0.51 0.415 0.51 0.56 0.385 0.56  ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 5.13 -0.085 5.13 0.085 4.875 0.085 4.875 0.235 4.74 0.235 4.74 0.085 4.13 0.085 4.13 0.42 3.995 0.42 3.995 0.085 2.895 0.085 2.895 0.21 2.76 0.21 2.76 0.085 1.9 0.085 1.9 0.32 1.83 0.32 1.83 0.085 1.55 0.085 1.55 0.21 1.415 0.21 1.415 0.085 1.135 0.085 1.135 0.285 1 0.285 1 0.085 0.34 0.085 0.34 0.32 0.27 0.32 0.27 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.375 0.92 0.93 0.92 0.93 0.485 1 0.485 1 0.99 0.51 0.99 0.51 1.12 0.375 1.12  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.365 0.56 1.46 0.56 1.46 0.7 1.365 0.7  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.085 0.29 0.155 0.29 0.155 0.785 0.865 0.785 0.865 0.855 0.18 0.855 0.18 1.145 0.085 1.145  ;
        POLYGON 1.225 0.25 1.36 0.25 1.36 0.415 1.63 0.415 1.63 0.485 1.295 0.485 1.295 0.795 1.325 0.795 1.325 0.93 1.225 0.93  ;
        POLYGON 0.65 1.055 1.065 1.055 1.065 0.42 0.625 0.42 0.625 0.325 0.76 0.325 0.76 0.35 1.135 0.35 1.135 1.055 1.295 1.055 1.295 1.18 1.695 1.18 1.695 1.25 1.225 1.25 1.225 1.125 0.65 1.125  ;
        POLYGON 1.65 0.795 1.695 0.795 1.695 0.35 1.635 0.35 1.635 0.215 1.765 0.215 1.765 0.645 2.11 0.645 2.11 0.715 1.765 0.715 1.765 0.93 1.65 0.93  ;
        POLYGON 2.065 0.45 2.245 0.45 2.245 0.9 2.175 0.9 2.175 0.52 2.065 0.52  ;
        POLYGON 2.445 0.525 2.955 0.525 2.955 0.44 3.09 0.44 3.09 0.645 3.175 0.645 3.175 0.715 3.02 0.715 3.02 0.595 2.445 0.595  ;
        POLYGON 2.14 0.965 2.31 0.965 2.31 0.305 2.175 0.305 2.175 0.235 2.38 0.235 2.38 0.965 2.95 0.965 2.95 0.78 3.22 0.78 3.22 0.765 3.355 0.765 3.355 0.85 3.02 0.85 3.02 1.035 2.21 1.035 2.21 1.185 2.14 1.185  ;
        POLYGON 3.375 0.41 3.445 0.41 3.445 0.545 3.66 0.545 3.66 0.895 3.59 0.895 3.59 0.615 3.375 0.615  ;
        POLYGON 3.515 0.96 3.725 0.96 3.725 0.48 3.51 0.48 3.51 0.41 3.795 0.41 3.795 0.78 4.37 0.78 4.37 0.85 3.795 0.85 3.795 1.03 3.515 1.03  ;
        POLYGON 3.86 0.915 4.45 0.915 4.45 0.51 4.405 0.51 4.405 0.235 4.52 0.235 4.52 0.985 3.86 0.985  ;
  END
END SDFFS_X2

MACRO SDFF_X1
  CLASS core ;
  FOREIGN SDFF_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 4.37 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.43 0.2 0.51 0.2 0.51 0.42 0.5 0.42 0.5 1.025 0.43 1.025  ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.67 0.765 3.865 0.765 3.865 0.98 3.67 0.98  ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.235 1.315 0.235 0.95 0.305 0.95 0.305 1.315 0.725 1.315 0.725 1.115 0.86 1.115 0.86 1.315 1.64 1.315 1.64 0.99 1.71 0.99 1.71 1.315 2.165 1.315 2.165 1.08 2.235 1.08 2.235 1.315 2.925 1.315 2.925 1.17 2.995 1.17 2.995 1.315 3.31 1.315 3.31 1.205 3.38 1.205 3.38 1.315 4.065 1.315 4.065 1.205 4.135 1.205 4.135 1.315 4.37 1.315 4.37 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.055 0.2 0.13 0.2 0.13 1.025 0.055 1.025  ;
    END
  END Q
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.385 0.915 3.48 0.915 3.48 0.63 4.06 0.63 4.06 0.7 3.55 0.7 3.55 0.985 3.385 0.985  ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 4.37 -0.085 4.37 0.085 4.14 0.085 4.14 0.195 4.07 0.195 4.07 0.085 3.415 0.085 3.415 0.16 3.28 0.16 3.28 0.085 2.995 0.085 2.995 0.28 2.925 0.28 2.925 0.085 2.235 0.085 2.235 0.37 2.165 0.37 2.165 0.085 1.705 0.085 1.705 0.445 1.635 0.445 1.635 0.085 0.955 0.085 0.955 0.41 0.82 0.41 0.82 0.085 0.31 0.085 0.31 0.32 0.24 0.32 0.24 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.99 0.77 4.125 0.77 4.125 0.565 3.42 0.565 3.42 0.37 3.49 0.37 3.49 0.495 4.195 0.495 4.195 1.02 3.99 1.02  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.015 0.7 3.17 0.7 3.17 0.84 3.015 0.84  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.565 1.075 0.585 1.075 0.585 0.185 0.73 0.185 0.73 0.46 0.655 0.46 0.655 1.21 0.565 1.21  ;
        POLYGON 0.72 0.915 0.795 0.915 0.795 0.475 1.08 0.475 1.08 0.36 1.36 0.36 1.36 0.43 1.15 0.43 1.15 0.545 0.865 0.545 0.865 0.98 1.205 0.98 1.205 1.2 1.135 1.2 1.135 1.05 0.72 1.05  ;
        POLYGON 1.02 0.845 1.335 0.845 1.335 0.605 1.825 0.605 1.825 0.415 1.895 0.415 1.895 1.02 1.825 1.02 1.825 0.675 1.405 0.675 1.405 0.915 1.02 0.915  ;
        POLYGON 1.96 0.25 2.05 0.25 2.05 0.56 2.3 0.56 2.3 0.695 2.05 0.695 2.05 1.2 1.96 1.2  ;
        POLYGON 2.435 1.115 2.65 1.115 2.65 1.185 2.365 1.185 2.365 0.975 2.115 0.975 2.115 0.84 2.365 0.84 2.365 0.27 2.65 0.27 2.65 0.34 2.435 0.34  ;
        POLYGON 2.57 0.98 3.185 0.98 3.185 1.115 3.115 1.115 3.115 1.05 2.5 1.05 2.5 0.405 3.115 0.405 3.115 0.25 3.185 0.25 3.185 0.475 2.57 0.475  ;
        POLYGON 3.32 1.05 3.79 1.05 3.79 1.12 3.25 1.12 3.25 0.635 2.815 0.635 2.815 0.565 3.25 0.565 3.25 0.225 3.655 0.225 3.655 0.2 3.79 0.2 3.79 0.295 3.32 0.295  ;
        POLYGON 3.575 0.36 4.26 0.36 4.26 0.165 4.335 0.165 4.335 1.145 4.26 1.145 4.26 0.43 3.575 0.43  ;
  END
END SDFF_X1

MACRO SDFF_X2
  CLASS core ;
  FOREIGN SDFF_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 4.37 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.425 0.28 0.51 0.28 0.51 0.42 0.495 0.42 0.495 1.25 0.425 1.25  ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.635 0.785 3.86 0.785 3.86 0.945 3.635 0.945  ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.205 1.315 0.205 1.065 0.34 1.065 0.34 1.315 0.745 1.315 0.745 1.115 0.88 1.115 0.88 1.315 1.52 1.315 1.52 1.115 1.655 1.115 1.655 1.315 2.11 1.315 2.11 1.115 2.245 1.115 2.245 1.315 2.87 1.315 2.87 1.115 3.005 1.115 3.005 1.315 3.24 1.315 3.24 1.205 3.375 1.205 3.375 1.315 4 1.315 4 1.065 4.135 1.065 4.135 1.315 4.37 1.315 4.37 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.05 0.28 0.13 0.28 0.13 1.11 0.05 1.11  ;
    END
  END Q
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.355 0.85 3.48 0.85 3.48 0.65 3.85 0.65 3.85 0.61 3.985 0.61 3.985 0.72 3.55 0.72 3.55 0.985 3.355 0.985  ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 4.37 -0.085 4.37 0.085 4.135 0.085 4.135 0.16 4 0.16 4 0.085 3.34 0.085 3.34 0.195 3.27 0.195 3.27 0.085 2.995 0.085 2.995 0.245 2.86 0.245 2.86 0.085 2.22 0.085 2.22 0.335 2.085 0.335 2.085 0.085 1.655 0.085 1.655 0.41 1.52 0.41 1.52 0.085 0.865 0.085 0.865 0.23 0.73 0.23 0.73 0.085 0.3 0.085 0.3 0.32 0.23 0.32 0.23 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.925 0.85 4.05 0.85 4.05 0.545 3.785 0.545 3.785 0.585 3.355 0.585 3.355 0.515 3.715 0.515 3.715 0.475 4.12 0.475 4.12 0.985 3.925 0.985  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.91 0.7 3.085 0.7 3.085 0.84 2.91 0.84  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.575 0.185 0.645 0.185 0.645 1.08 0.66 1.08 0.66 1.215 0.575 1.215  ;
        POLYGON 0.78 0.955 1.28 0.955 1.28 1.025 0.71 1.025 0.71 0.36 1.26 0.36 1.26 0.43 0.78 0.43  ;
        POLYGON 1.045 0.795 1.71 0.795 1.71 0.565 1.29 0.565 1.29 0.495 1.71 0.495 1.71 0.45 1.845 0.45 1.845 1.075 1.71 1.075 1.71 0.865 1.045 0.865  ;
        POLYGON 1.91 0.25 1.99 0.25 1.99 0.91 2.28 0.91 2.28 1.045 2.045 1.045 2.045 1.165 1.91 1.165  ;
        POLYGON 2.415 1.095 2.62 1.095 2.62 1.165 2.345 1.165 2.345 0.555 2.055 0.555 2.055 0.42 2.345 0.42 2.345 0.285 2.6 0.285 2.6 0.355 2.415 0.355  ;
        POLYGON 2.735 0.935 3.155 0.935 3.155 1.11 3.085 1.11 3.085 1.005 2.48 1.005 2.48 0.85 2.665 0.85 2.665 0.315 3.08 0.315 3.08 0.25 3.15 0.25 3.15 0.385 2.735 0.385  ;
        POLYGON 3.29 1.05 3.75 1.05 3.75 1.12 3.22 1.12 3.22 0.635 2.8 0.635 2.8 0.565 3.22 0.565 3.22 0.345 3.405 0.345 3.405 0.165 3.75 0.165 3.75 0.235 3.475 0.235 3.475 0.415 3.29 0.415  ;
        POLYGON 3.545 0.305 4.215 0.305 4.215 0.165 4.285 0.165 4.285 1.25 4.215 1.25 4.215 0.375 3.615 0.375 3.615 0.44 3.545 0.44  ;
  END
END SDFF_X2

MACRO TBUF_X1
  CLASS core ;
  FOREIGN TBUF_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.205 0.71 0.205 0.71 0.275 0.51 0.275 0.51 1 0.675 1 0.675 1.22 0.605 1.22 0.605 1.07 0.44 1.07  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.17 0.56 0.32 0.56 0.32 0.7 0.17 0.7  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.225 1.315 0.225 1.145 0.295 1.145 0.295 1.315 0.755 1.315 0.755 0.86 0.825 0.86 0.825 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 1.06 0.085 1.06 0.23 0.99 0.23 0.99 0.085 0.295 0.085 0.295 0.265 0.225 0.265 0.225 0.085 0 0.085  ;
    END
  END VSS
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.785 0.53 0.98 0.53 0.98 0.665 0.785 0.665  ;
    END
  END EN
  OBS
      LAYER metal1 ;
        POLYGON 0.035 0.15 0.11 0.15 0.11 0.425 0.375 0.425 0.375 0.495 0.105 0.495 0.105 1.085 0.11 1.085 0.11 1.22 0.035 1.22  ;
        POLYGON 0.575 0.34 0.775 0.34 0.775 0.15 0.91 0.15 0.91 0.41 0.645 0.41 0.645 0.935 0.575 0.935  ;
  END
END TBUF_X1

MACRO TBUF_X16
  CLASS core ;
  FOREIGN TBUF_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 3.61 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.54 0.265 3.01 0.265 3.01 0.335 0.61 0.335 0.61 0.7 2.98 0.7 2.98 1.04 2.91 1.04 2.91 0.77 2.22 0.77 2.22 1.04 2.15 1.04 2.15 0.77 1.46 0.77 1.46 1.04 1.39 1.04 1.39 0.77 0.7 0.77 0.7 1.04 0.54 1.04  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2 0.425 0.355 0.425 0.355 0.525 0.27 0.525 0.27 0.56 0.2 0.56  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.245 1.315 0.245 1.08 0.315 1.08 0.315 1.315 1.005 1.315 1.005 0.94 1.075 0.94 1.075 1.315 1.765 1.315 1.765 0.94 1.835 0.94 1.835 1.315 2.525 1.315 2.525 0.94 2.595 0.94 2.595 1.315 3.285 1.315 3.285 0.82 3.355 0.82 3.355 1.315 3.61 1.315 3.61 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 3.61 -0.085 3.61 0.085 3.36 0.085 3.36 0.265 3.29 0.265 3.29 0.085 2.595 0.085 2.595 0.195 2.525 0.195 2.525 0.085 1.835 0.085 1.835 0.195 1.765 0.195 1.765 0.085 1.075 0.085 1.075 0.195 1.005 0.195 1.005 0.085 0.315 0.085 0.315 0.36 0.245 0.36 0.245 0.085 0 0.085  ;
    END
  END VSS
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.29 0.56 3.415 0.56 3.415 0.7 3.29 0.7  ;
    END
  END EN
  OBS
      LAYER metal1 ;
        POLYGON 0.035 0.245 0.13 0.245 0.13 0.67 0.335 0.67 0.335 0.595 0.47 0.595 0.47 0.74 0.13 0.74 0.13 1.155 0.035 1.155  ;
        POLYGON 0.675 0.4 3.48 0.4 3.48 0.15 3.575 0.15 3.575 0.9 3.48 0.9 3.48 0.47 0.675 0.47  ;
  END
END TBUF_X16

MACRO TBUF_X2
  CLASS core ;
  FOREIGN TBUF_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.51 0.69 0.675 0.69 0.675 1.165 0.605 1.165 0.605 0.76 0.44 0.76 0.44 0.355 0.605 0.355 0.605 0.15 0.675 0.15 0.675 0.425 0.51 0.425  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.215 0.56 0.215 0.7 0.06 0.7  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.225 1.315 0.225 1.175 0.295 1.175 0.295 1.315 0.945 1.315 0.945 1.175 1.015 1.175 1.015 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 1.02 0.085 1.02 0.265 0.95 0.265 0.95 0.085 0.295 0.085 0.295 0.265 0.225 0.265 0.225 0.085 0 0.085  ;
    END
  END VSS
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.875 0.7 1.08 0.7 1.08 0.875 0.875 0.875  ;
    END
  END EN
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.765 0.305 0.765 0.305 0.4 0.045 0.4 0.045 0.15 0.115 0.15 0.115 0.33 0.375 0.33 0.375 0.835 0.115 0.835 0.115 1.25 0.045 1.25  ;
        POLYGON 0.575 0.49 0.74 0.49 0.74 0.15 0.835 0.15 0.835 0.285 0.81 0.285 0.81 1.115 0.83 1.115 0.83 1.25 0.74 1.25 0.74 0.625 0.575 0.625  ;
  END
END TBUF_X2

MACRO TBUF_X4
  CLASS core ;
  FOREIGN TBUF_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.33 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.615 0.765 0.7 0.765 0.7 1.04 0.545 1.04 0.545 0.205 0.695 0.205 0.695 0.34 0.615 0.34  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.19 0.56 0.32 0.56 0.32 0.7 0.19 0.7  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.245 1.315 0.245 1.08 0.315 1.08 0.315 1.315 1.005 1.315 1.005 0.82 1.075 0.82 1.075 1.315 1.33 1.315 1.33 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.33 -0.085 1.33 0.085 1.08 0.085 1.08 0.265 1.01 0.265 1.01 0.085 0.315 0.085 0.315 0.36 0.245 0.36 0.245 0.085 0 0.085  ;
    END
  END VSS
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.01 0.56 1.135 0.56 1.135 0.7 1.01 0.7  ;
    END
  END EN
  OBS
      LAYER metal1 ;
        POLYGON 0.055 0.245 0.13 0.245 0.13 0.425 0.455 0.425 0.455 0.655 0.385 0.655 0.385 0.495 0.125 0.495 0.125 1.02 0.13 1.02 0.13 1.155 0.055 1.155  ;
        POLYGON 0.68 0.405 1.2 0.405 1.2 0.15 1.295 0.15 1.295 0.9 1.2 0.9 1.2 0.475 0.68 0.475  ;
  END
END TBUF_X4

MACRO TBUF_X8
  CLASS core ;
  FOREIGN TBUF_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.09 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.54 0.235 1.46 0.235 1.46 1.04 1.39 1.04 1.39 0.305 0.61 0.305 0.61 0.835 0.7 0.835 0.7 1.11 0.54 1.11  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.175 0.56 0.32 0.56 0.32 0.7 0.175 0.7  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.25 1.315 0.25 1.08 0.32 1.08 0.32 1.315 1.01 1.315 1.01 0.94 1.08 0.94 1.08 1.315 1.77 1.315 1.77 1.08 1.84 1.08 1.84 1.315 2.09 1.315 2.09 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.09 -0.085 2.09 0.085 1.845 0.085 1.845 0.36 1.775 0.36 1.775 0.085 1.12 0.085 1.12 0.16 0.985 0.16 0.985 0.085 0.32 0.085 0.32 0.36 0.25 0.36 0.25 0.085 0 0.085  ;
    END
  END VSS
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.685 0.67 1.255 0.67 1.255 0.635 1.325 0.635 1.325 0.77 0.685 0.77  ;
        POLYGON 1.525 0.635 1.92 0.635 1.92 0.705 1.65 0.705 1.65 0.84 1.525 0.84  ;
    END
  END EN
  OBS
      LAYER metal1 ;
        POLYGON 0.04 0.245 0.135 0.245 0.135 0.425 0.455 0.425 0.455 0.56 0.385 0.56 0.385 0.495 0.11 0.495 0.11 1.02 0.135 1.02 0.135 1.155 0.04 1.155  ;
        POLYGON 0.675 0.405 1.255 0.405 1.255 0.37 1.325 0.37 1.325 0.505 0.675 0.505  ;
        POLYGON 1.965 1.02 1.985 1.02 1.985 0.505 1.525 0.505 1.525 0.37 1.595 0.37 1.595 0.435 1.965 0.435 1.965 0.245 2.055 0.245 2.055 1.155 1.965 1.155  ;
  END
END TBUF_X8

MACRO TINV_X1
  CLASS core ;
  FOREIGN TINV_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.225 1.315 0.225 1.145 0.295 1.145 0.295 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.295 0.085 0.295 0.295 0.225 0.295 0.225 0.085 0 0.085  ;
    END
  END VSS
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.215 0.595 0.385 0.595 0.385 0.665 0.215 0.665  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.61 1.105 0.655 1.105 0.655 0.275 0.405 0.275 0.405 0.175 0.725 0.175 0.725 1.24 0.61 1.24  ;
    END
  END ZN
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.17 0.945 0.44 0.945 0.44 0.7 0.55 0.7 0.55 1.08 0.17 1.08  ;
    END
  END EN
  OBS
      LAYER metal1 ;
        POLYGON 0.035 0.175 0.11 0.175 0.11 0.375 0.59 0.375 0.59 0.445 0.105 0.445 0.105 1.105 0.11 1.105 0.11 1.24 0.035 1.24  ;
  END
END TINV_X1

MACRO TLAT_X1
  CLASS core ;
  FOREIGN TLAT_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.47 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.3 1.315 0.3 0.885 0.37 0.885 0.37 1.315 0.645 1.315 0.645 0.94 0.715 0.94 0.715 1.315 1.38 1.315 1.38 1.115 1.515 1.115 1.515 1.315 2.365 1.315 2.365 1.115 1.93 1.115 1.93 1 2.065 1 2.065 1.045 2.435 1.045 2.435 1.315 2.47 1.315 2.47 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.34 0.28 2.41 0.28 2.41 0.98 2.34 0.98  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.47 -0.085 2.47 0.085 2.025 0.085 2.025 0.45 1.955 0.45 1.955 0.085 1.47 0.085 1.47 0.32 1.4 0.32 1.4 0.085 0.72 0.085 0.72 0.32 0.65 0.32 0.65 0.085 0.37 0.085 0.37 0.245 0.3 0.245 0.3 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.73 0.42 0.89 0.42 0.89 0.56 0.73 0.56  ;
    END
  END D
  PIN OE
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.39 0.84 1.56 0.84 1.56 1.035 1.39 1.035  ;
    END
  END OE
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2 0.56 0.32 0.56 0.32 0.7 0.2 0.7  ;
    END
  END G
  OBS
      LAYER metal1 ;
        POLYGON 0.065 0.215 0.185 0.215 0.185 0.37 0.43 0.37 0.43 0.505 0.36 0.505 0.36 0.44 0.135 0.44 0.135 0.765 0.185 0.765 0.185 1.04 0.065 1.04  ;
        POLYGON 0.495 0.215 0.585 0.215 0.585 0.805 0.95 0.805 0.95 0.59 1.02 0.59 1.02 0.875 0.495 0.875  ;
        POLYGON 1.595 0.185 1.705 0.185 1.705 0.46 1.595 0.46  ;
        POLYGON 1.03 0.94 1.085 0.94 1.085 0.395 0.995 0.395 0.995 0.325 1.155 0.325 1.155 0.66 1.955 0.66 1.955 0.73 1.155 0.73 1.155 1.215 1.03 1.215  ;
        POLYGON 1.775 0.865 2.02 0.865 2.02 0.595 1.29 0.595 1.29 0.525 1.77 0.525 1.77 0.42 1.84 0.42 1.84 0.525 2.09 0.525 2.09 0.935 1.845 0.935 1.845 1.025 1.775 1.025  ;
        POLYGON 1.6 1.115 1.635 1.115 1.635 0.795 1.705 0.795 1.705 1.18 2.3 1.18 2.3 1.25 1.6 1.25  ;
  END
END TLAT_X1

MACRO XNOR2_X1
  CLASS core ;
  FOREIGN XNOR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.175 0.42 0.32 0.42 0.32 0.49 0.755 0.49 0.755 0.56 0.175 0.56  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.145 0.11 1.145 0.11 1.315 0.42 1.315 0.42 1.145 0.49 1.145 0.49 1.315 1 1.315 1 1.205 1.07 1.205 1.07 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.49 0.085 0.49 0.365 0.42 0.365 0.42 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.36 0.845 0.43 0.845 0.43 0.91 0.63 0.91 0.63 0.84 0.97 0.84 0.97 0.98 0.36 0.98  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 1.045 1.035 1.045 1.035 0.56 0.82 0.56 0.82 0.285 0.89 0.285 0.89 0.49 1.105 0.49 1.105 1.115 0.7 1.115 0.7 1.22 0.63 1.22  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.04 0.285 0.11 0.285 0.11 0.71 0.565 0.71 0.565 0.845 0.495 0.845 0.495 0.78 0.295 0.78 0.295 1.22 0.225 1.22 0.225 0.78 0.04 0.78  ;
        POLYGON 0.63 0.15 1.07 0.15 1.07 0.365 1 0.365 1 0.22 0.7 0.22 0.7 0.365 0.63 0.365  ;
  END
END XNOR2_X1

MACRO XNOR2_X2
  CLASS core ;
  FOREIGN XNOR2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.17 0.49 0.44 0.49 0.44 0.42 0.51 0.42 0.51 0.49 0.825 0.49 0.825 0.56 0.17 0.56  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.055 1.315 0.055 1.17 0.125 1.17 0.125 1.315 0.43 1.315 0.43 1.17 0.5 1.17 0.5 1.315 1.015 1.315 1.015 1.17 1.085 1.17 1.085 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.52 0.085 0.52 0.24 0.45 0.24 0.45 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.32 0.695 0.945 0.695 0.945 0.84 0.82 0.84 0.82 0.765 0.32 0.765  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.645 0.975 1.01 0.975 1.01 0.42 0.8 0.42 0.8 0.325 0.935 0.325 0.935 0.35 1.08 0.35 1.08 1.045 0.715 1.045 0.715 1.25 0.645 1.25  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.105 0.83 0.58 0.83 0.58 0.905 0.31 0.905 0.31 1.245 0.24 1.245 0.24 0.905 0.035 0.905 0.035 0.29 0.125 0.29 0.125 0.425 0.105 0.425  ;
        POLYGON 0.645 0.15 1.085 0.15 1.085 0.285 1.015 0.285 1.015 0.22 0.715 0.22 0.715 0.285 0.645 0.285  ;
  END
END XNOR2_X2

MACRO XOR2_X1
  CLASS core ;
  FOREIGN XOR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.805 0.965 1.035 0.965 1.035 0.42 0.63 0.42 0.63 0.285 0.615 0.285 0.615 0.15 0.7 0.15 0.7 0.35 1.105 0.35 1.105 1.035 0.875 1.035 0.875 1.115 0.805 1.115  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.175 0.84 0.74 0.84 0.74 0.98 0.175 0.98  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.42 1.315 0.42 1.1 0.49 1.1 0.49 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 1.055 0.085 1.055 0.27 0.985 0.27 0.985 0.085 0.49 0.085 0.49 0.27 0.42 0.27 0.42 0.085 0.11 0.085 0.11 0.27 0.04 0.27 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.34 0.56 0.97 0.56 0.97 0.7 0.34 0.7  ;
    END
  END B
  OBS
      LAYER metal1 ;
        POLYGON 0.04 0.34 0.225 0.34 0.225 0.15 0.295 0.15 0.295 0.34 0.565 0.34 0.565 0.425 0.11 0.425 0.11 1.115 0.04 1.115  ;
        POLYGON 0.615 1.1 0.685 1.1 0.685 1.18 0.985 1.18 0.985 1.1 1.055 1.1 1.055 1.25 0.615 1.25  ;
  END
END XOR2_X1

MACRO XOR2_X2
  CLASS core ;
  FOREIGN XOR2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.82 0.765 1.035 0.765 1.035 0.42 0.595 0.42 0.595 0.28 1.105 0.28 1.105 0.835 0.89 0.835 0.89 1.025 0.82 1.025  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.175 0.795 0.755 0.795 0.755 0.865 0.32 0.865 0.32 0.98 0.175 0.98  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.42 1.315 0.42 1.205 0.49 1.205 0.49 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 1.07 0.085 1.07 0.195 1 0.195 1 0.085 0.485 0.085 0.485 0.275 0.415 0.275 0.415 0.085 0.11 0.085 0.11 0.275 0.04 0.275 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.56 0.38 0.56 0.38 0.625 0.97 0.625 0.97 0.7 0.25 0.7  ;
    END
  END B
  OBS
      LAYER metal1 ;
        POLYGON 0.035 0.37 0.225 0.37 0.225 0.155 0.295 0.155 0.295 0.37 0.53 0.37 0.53 0.505 0.46 0.505 0.46 0.44 0.11 0.44 0.11 1.22 0.035 1.22  ;
        POLYGON 0.595 1.125 1.105 1.125 1.105 1.195 0.595 1.195  ;
  END
END XOR2_X2

END LIBRARY
#
# End of file
#
